
module ahb_slave_ram ( clk, reset, HSEL, HADDR, HBURST, HSIZE, HTRANS, HWRITE, 
        HWDATA, RANDSPLIT, HMASTER, HMASTLOCK, HRDATA, HREADY, HRESP, HSPLIT, 
        WR, RD, ADDR_WR, ADDR_RD, DIN, DOUT, STALL_pre );
  input [23:0] HADDR;
  input [2:0] HBURST;
  input [1:0] HSIZE;
  input [1:0] HTRANS;
  input [31:0] HWDATA;
  input [2:0] RANDSPLIT;
  input [3:0] HMASTER;
  output [31:0] HRDATA;
  output [1:0] HRESP;
  output [15:0] HSPLIT;
  output [8:0] ADDR_WR;
  output [8:0] ADDR_RD;
  output [31:0] DIN;
  input [31:0] DOUT;
  input clk, reset, HSEL, HWRITE, HMASTLOCK, STALL_pre;
  output HREADY, WR, RD;
  wire   STALL, split, N34, N35, N36, N37, N56, N57, data_phase, WR_pre_d, n68,
         n69, n71, n72, n73, n74, n75, n76, n77, n78, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n126, n127, n128, n129, n131, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n2, n3, n39, n40, n41, n42, n44, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70;
  wire   [2:0] waitstate;
  wire   [2:0] waitstate_pre;

  DFFSR STALL_reg ( .D(STALL_pre), .CLK(clk), .R(n52), .S(1'b1), .Q(STALL) );
  AND2X2 U42 ( .A(HMASTER[0]), .B(n101), .Y(n84) );
  AND2X2 U43 ( .A(n101), .B(n70), .Y(n87) );
  AND2X2 U44 ( .A(HMASTER[3]), .B(n104), .Y(n101) );
  AND2X2 U45 ( .A(n121), .B(HMASTER[0]), .Y(n107) );
  AND2X2 U46 ( .A(n121), .B(n70), .Y(n110) );
  AND2X2 U47 ( .A(RANDSPLIT[1]), .B(split), .Y(N57) );
  AND2X2 U48 ( .A(RANDSPLIT[0]), .B(split), .Y(N56) );
  AND2X2 U49 ( .A(n140), .B(n141), .Y(n139) );
  AND2X2 U50 ( .A(DOUT[9]), .B(n44), .Y(HRDATA[9]) );
  AND2X2 U51 ( .A(DOUT[8]), .B(n44), .Y(HRDATA[8]) );
  AND2X2 U52 ( .A(DOUT[7]), .B(n44), .Y(HRDATA[7]) );
  AND2X2 U53 ( .A(DOUT[6]), .B(n44), .Y(HRDATA[6]) );
  AND2X2 U54 ( .A(DOUT[5]), .B(n44), .Y(HRDATA[5]) );
  AND2X2 U55 ( .A(DOUT[4]), .B(n44), .Y(HRDATA[4]) );
  AND2X2 U56 ( .A(DOUT[3]), .B(n44), .Y(HRDATA[3]) );
  AND2X2 U57 ( .A(DOUT[31]), .B(n44), .Y(HRDATA[31]) );
  AND2X2 U58 ( .A(DOUT[30]), .B(n44), .Y(HRDATA[30]) );
  AND2X2 U59 ( .A(DOUT[2]), .B(n44), .Y(HRDATA[2]) );
  AND2X2 U60 ( .A(DOUT[29]), .B(n44), .Y(HRDATA[29]) );
  AND2X2 U61 ( .A(DOUT[28]), .B(n44), .Y(HRDATA[28]) );
  AND2X2 U62 ( .A(DOUT[27]), .B(n44), .Y(HRDATA[27]) );
  AND2X2 U63 ( .A(DOUT[26]), .B(n44), .Y(HRDATA[26]) );
  AND2X2 U64 ( .A(DOUT[25]), .B(n44), .Y(HRDATA[25]) );
  AND2X2 U65 ( .A(DOUT[24]), .B(n44), .Y(HRDATA[24]) );
  AND2X2 U66 ( .A(DOUT[23]), .B(n44), .Y(HRDATA[23]) );
  AND2X2 U67 ( .A(DOUT[22]), .B(n44), .Y(HRDATA[22]) );
  AND2X2 U68 ( .A(DOUT[21]), .B(n44), .Y(HRDATA[21]) );
  AND2X2 U69 ( .A(DOUT[20]), .B(n44), .Y(HRDATA[20]) );
  AND2X2 U70 ( .A(DOUT[1]), .B(n44), .Y(HRDATA[1]) );
  AND2X2 U71 ( .A(DOUT[19]), .B(n44), .Y(HRDATA[19]) );
  AND2X2 U72 ( .A(DOUT[18]), .B(n44), .Y(HRDATA[18]) );
  AND2X2 U73 ( .A(DOUT[17]), .B(n44), .Y(HRDATA[17]) );
  AND2X2 U74 ( .A(DOUT[16]), .B(n44), .Y(HRDATA[16]) );
  AND2X2 U75 ( .A(DOUT[15]), .B(n44), .Y(HRDATA[15]) );
  AND2X2 U76 ( .A(DOUT[14]), .B(n44), .Y(HRDATA[14]) );
  AND2X2 U77 ( .A(DOUT[13]), .B(n44), .Y(HRDATA[13]) );
  AND2X2 U78 ( .A(DOUT[12]), .B(n44), .Y(HRDATA[12]) );
  AND2X2 U79 ( .A(DOUT[11]), .B(n44), .Y(HRDATA[11]) );
  AND2X2 U80 ( .A(DOUT[10]), .B(n44), .Y(HRDATA[10]) );
  AND2X2 U81 ( .A(DOUT[0]), .B(n44), .Y(HRDATA[0]) );
  AND2X2 U82 ( .A(HWDATA[9]), .B(HREADY), .Y(DIN[9]) );
  AND2X2 U83 ( .A(HWDATA[8]), .B(HREADY), .Y(DIN[8]) );
  AND2X2 U84 ( .A(HWDATA[7]), .B(HREADY), .Y(DIN[7]) );
  AND2X2 U85 ( .A(HWDATA[6]), .B(HREADY), .Y(DIN[6]) );
  AND2X2 U86 ( .A(HWDATA[5]), .B(HREADY), .Y(DIN[5]) );
  AND2X2 U87 ( .A(HWDATA[4]), .B(HREADY), .Y(DIN[4]) );
  AND2X2 U88 ( .A(HWDATA[3]), .B(HREADY), .Y(DIN[3]) );
  AND2X2 U89 ( .A(HWDATA[31]), .B(HREADY), .Y(DIN[31]) );
  AND2X2 U90 ( .A(HWDATA[30]), .B(HREADY), .Y(DIN[30]) );
  AND2X2 U91 ( .A(HWDATA[2]), .B(HREADY), .Y(DIN[2]) );
  AND2X2 U92 ( .A(HWDATA[29]), .B(HREADY), .Y(DIN[29]) );
  AND2X2 U93 ( .A(HWDATA[28]), .B(HREADY), .Y(DIN[28]) );
  AND2X2 U94 ( .A(HWDATA[27]), .B(HREADY), .Y(DIN[27]) );
  AND2X2 U95 ( .A(HWDATA[26]), .B(HREADY), .Y(DIN[26]) );
  AND2X2 U96 ( .A(HWDATA[25]), .B(HREADY), .Y(DIN[25]) );
  AND2X2 U97 ( .A(HWDATA[24]), .B(HREADY), .Y(DIN[24]) );
  AND2X2 U98 ( .A(HWDATA[23]), .B(HREADY), .Y(DIN[23]) );
  AND2X2 U99 ( .A(HWDATA[22]), .B(HREADY), .Y(DIN[22]) );
  AND2X2 U100 ( .A(HWDATA[21]), .B(HREADY), .Y(DIN[21]) );
  AND2X2 U101 ( .A(HWDATA[20]), .B(HREADY), .Y(DIN[20]) );
  AND2X2 U102 ( .A(HWDATA[1]), .B(HREADY), .Y(DIN[1]) );
  AND2X2 U103 ( .A(HWDATA[19]), .B(HREADY), .Y(DIN[19]) );
  AND2X2 U104 ( .A(HWDATA[18]), .B(HREADY), .Y(DIN[18]) );
  AND2X2 U105 ( .A(HWDATA[17]), .B(HREADY), .Y(DIN[17]) );
  AND2X2 U106 ( .A(HWDATA[16]), .B(HREADY), .Y(DIN[16]) );
  AND2X2 U107 ( .A(HWDATA[15]), .B(HREADY), .Y(DIN[15]) );
  AND2X2 U108 ( .A(HWDATA[14]), .B(HREADY), .Y(DIN[14]) );
  AND2X2 U109 ( .A(HWDATA[13]), .B(HREADY), .Y(DIN[13]) );
  AND2X2 U110 ( .A(HWDATA[12]), .B(HREADY), .Y(DIN[12]) );
  AND2X2 U111 ( .A(HWDATA[11]), .B(HREADY), .Y(DIN[11]) );
  AND2X2 U112 ( .A(HWDATA[10]), .B(HREADY), .Y(DIN[10]) );
  AND2X2 U113 ( .A(HWDATA[0]), .B(HREADY), .Y(DIN[0]) );
  OAI21X1 U137 ( .A(HREADY), .B(n51), .C(n68), .Y(n154) );
  OAI21X1 U138 ( .A(n68), .B(n62), .C(n69), .Y(n155) );
  NAND2X1 U139 ( .A(ADDR_WR[0]), .B(n46), .Y(n69) );
  OAI21X1 U140 ( .A(n68), .B(n61), .C(n71), .Y(n156) );
  NAND2X1 U141 ( .A(ADDR_WR[1]), .B(n46), .Y(n71) );
  OAI21X1 U142 ( .A(n68), .B(n60), .C(n72), .Y(n157) );
  NAND2X1 U143 ( .A(ADDR_WR[2]), .B(n46), .Y(n72) );
  OAI21X1 U144 ( .A(n68), .B(n59), .C(n73), .Y(n158) );
  NAND2X1 U145 ( .A(ADDR_WR[3]), .B(n46), .Y(n73) );
  OAI21X1 U146 ( .A(n68), .B(n58), .C(n74), .Y(n159) );
  NAND2X1 U147 ( .A(ADDR_WR[4]), .B(n46), .Y(n74) );
  OAI21X1 U148 ( .A(n68), .B(n57), .C(n75), .Y(n160) );
  NAND2X1 U149 ( .A(ADDR_WR[5]), .B(n46), .Y(n75) );
  OAI21X1 U150 ( .A(n68), .B(n56), .C(n76), .Y(n161) );
  NAND2X1 U151 ( .A(ADDR_WR[6]), .B(n46), .Y(n76) );
  OAI21X1 U152 ( .A(n68), .B(n55), .C(n77), .Y(n162) );
  NAND2X1 U153 ( .A(ADDR_WR[7]), .B(n46), .Y(n77) );
  OAI21X1 U154 ( .A(n68), .B(n54), .C(n78), .Y(n163) );
  NAND2X1 U155 ( .A(ADDR_WR[8]), .B(n46), .Y(n78) );
  NAND3X1 U156 ( .A(HTRANS[1]), .B(HREADY), .C(HWRITE), .Y(n68) );
  OAI21X1 U157 ( .A(HREADY), .B(n50), .C(n40), .Y(n164) );
  OAI21X1 U158 ( .A(n80), .B(n41), .C(n82), .Y(n165) );
  NAND2X1 U159 ( .A(HSPLIT[15]), .B(n80), .Y(n82) );
  NAND2X1 U160 ( .A(n83), .B(n84), .Y(n80) );
  OAI21X1 U161 ( .A(n42), .B(n85), .C(n86), .Y(n166) );
  NAND2X1 U162 ( .A(HSPLIT[14]), .B(n85), .Y(n86) );
  NAND2X1 U163 ( .A(n87), .B(n83), .Y(n85) );
  OAI21X1 U164 ( .A(n42), .B(n88), .C(n89), .Y(n167) );
  NAND2X1 U165 ( .A(HSPLIT[13]), .B(n88), .Y(n89) );
  NAND2X1 U166 ( .A(n90), .B(n84), .Y(n88) );
  OAI21X1 U167 ( .A(n41), .B(n91), .C(n92), .Y(n168) );
  NAND2X1 U168 ( .A(HSPLIT[12]), .B(n91), .Y(n92) );
  NAND2X1 U169 ( .A(n90), .B(n87), .Y(n91) );
  OAI21X1 U170 ( .A(n41), .B(n93), .C(n94), .Y(n169) );
  NAND2X1 U171 ( .A(HSPLIT[11]), .B(n93), .Y(n94) );
  NAND2X1 U172 ( .A(n95), .B(n84), .Y(n93) );
  OAI21X1 U173 ( .A(n42), .B(n96), .C(n97), .Y(n170) );
  NAND2X1 U174 ( .A(HSPLIT[10]), .B(n96), .Y(n97) );
  NAND2X1 U175 ( .A(n95), .B(n87), .Y(n96) );
  OAI21X1 U176 ( .A(n42), .B(n98), .C(n99), .Y(n171) );
  NAND2X1 U177 ( .A(HSPLIT[9]), .B(n98), .Y(n99) );
  NAND2X1 U178 ( .A(n100), .B(n84), .Y(n98) );
  OAI21X1 U179 ( .A(n41), .B(n102), .C(n103), .Y(n172) );
  NAND2X1 U180 ( .A(HSPLIT[8]), .B(n102), .Y(n103) );
  NAND2X1 U181 ( .A(n100), .B(n87), .Y(n102) );
  OAI21X1 U182 ( .A(n41), .B(n105), .C(n106), .Y(n173) );
  NAND2X1 U183 ( .A(HSPLIT[7]), .B(n105), .Y(n106) );
  NAND2X1 U184 ( .A(n107), .B(n83), .Y(n105) );
  OAI21X1 U185 ( .A(n42), .B(n108), .C(n109), .Y(n174) );
  NAND2X1 U186 ( .A(HSPLIT[6]), .B(n108), .Y(n109) );
  NAND2X1 U187 ( .A(n110), .B(n83), .Y(n108) );
  NOR2X1 U188 ( .A(n66), .B(n67), .Y(n83) );
  OAI21X1 U189 ( .A(n42), .B(n111), .C(n112), .Y(n175) );
  NAND2X1 U190 ( .A(HSPLIT[5]), .B(n111), .Y(n112) );
  NAND2X1 U191 ( .A(n107), .B(n90), .Y(n111) );
  OAI21X1 U192 ( .A(n41), .B(n113), .C(n114), .Y(n176) );
  NAND2X1 U193 ( .A(HSPLIT[4]), .B(n113), .Y(n114) );
  NAND2X1 U194 ( .A(n110), .B(n90), .Y(n113) );
  NOR2X1 U195 ( .A(n66), .B(HMASTER[1]), .Y(n90) );
  OAI21X1 U196 ( .A(n41), .B(n115), .C(n116), .Y(n177) );
  NAND2X1 U197 ( .A(HSPLIT[3]), .B(n115), .Y(n116) );
  NAND2X1 U198 ( .A(n107), .B(n95), .Y(n115) );
  OAI21X1 U199 ( .A(n42), .B(n117), .C(n118), .Y(n178) );
  NAND2X1 U200 ( .A(HSPLIT[2]), .B(n117), .Y(n118) );
  NAND2X1 U201 ( .A(n110), .B(n95), .Y(n117) );
  NOR2X1 U202 ( .A(n67), .B(HMASTER[2]), .Y(n95) );
  OAI21X1 U203 ( .A(n42), .B(n119), .C(n120), .Y(n179) );
  NAND2X1 U204 ( .A(HSPLIT[1]), .B(n119), .Y(n120) );
  NAND2X1 U205 ( .A(n107), .B(n100), .Y(n119) );
  OAI21X1 U206 ( .A(n41), .B(n122), .C(n123), .Y(n180) );
  NAND2X1 U207 ( .A(HSPLIT[0]), .B(n122), .Y(n123) );
  NAND2X1 U208 ( .A(n110), .B(n100), .Y(n122) );
  NOR2X1 U209 ( .A(HMASTER[1]), .B(HMASTER[2]), .Y(n100) );
  NOR2X1 U210 ( .A(n53), .B(HMASTER[3]), .Y(n121) );
  OAI21X1 U211 ( .A(split), .B(n65), .C(n124), .Y(n181) );
  OAI21X1 U212 ( .A(n3), .B(n126), .C(split), .Y(n124) );
  NAND2X1 U213 ( .A(n127), .B(n128), .Y(n126) );
  XOR2X1 U214 ( .A(n129), .B(waitstate[2]), .Y(n128) );
  XOR2X1 U216 ( .A(n48), .B(n131), .Y(n127) );
  XOR2X1 U217 ( .A(waitstate_pre[1]), .B(waitstate_pre[0]), .Y(n131) );
  NAND2X1 U220 ( .A(waitstate_pre[1]), .B(waitstate_pre[0]), .Y(n129) );
  NOR2X1 U221 ( .A(n51), .B(n46), .Y(WR) );
  OAI21X1 U222 ( .A(n133), .B(n49), .C(n134), .Y(N37) );
  NAND3X1 U223 ( .A(waitstate[1]), .B(waitstate[0]), .C(n135), .Y(n134) );
  NOR2X1 U224 ( .A(waitstate[2]), .B(n41), .Y(n135) );
  AOI21X1 U225 ( .A(n47), .B(n48), .C(N35), .Y(n133) );
  NOR2X1 U226 ( .A(n136), .B(n42), .Y(N36) );
  XOR2X1 U227 ( .A(waitstate[0]), .B(n48), .Y(n136) );
  NOR2X1 U228 ( .A(n42), .B(waitstate[0]), .Y(N35) );
  NAND2X1 U229 ( .A(n41), .B(n104), .Y(N34) );
  NAND2X1 U230 ( .A(split), .B(n104), .Y(n81) );
  NAND3X1 U231 ( .A(n137), .B(n138), .C(n139), .Y(n104) );
  NOR2X1 U232 ( .A(n142), .B(n143), .Y(n141) );
  NAND3X1 U233 ( .A(HADDR[17]), .B(HADDR[16]), .C(HADDR[18]), .Y(n143) );
  NAND3X1 U234 ( .A(HADDR[14]), .B(HADDR[13]), .C(HADDR[15]), .Y(n142) );
  NOR2X1 U235 ( .A(n144), .B(n145), .Y(n140) );
  NAND3X1 U236 ( .A(HADDR[23]), .B(HADDR[22]), .C(HADDR[9]), .Y(n145) );
  NAND3X1 U237 ( .A(HADDR[20]), .B(HADDR[19]), .C(HADDR[21]), .Y(n144) );
  NOR2X1 U238 ( .A(n146), .B(n147), .Y(n138) );
  NAND3X1 U239 ( .A(HADDR[4]), .B(HADDR[3]), .C(HADDR[5]), .Y(n147) );
  NAND3X1 U240 ( .A(HADDR[2]), .B(HADDR[1]), .C(n63), .Y(n146) );
  OAI21X1 U241 ( .A(HTRANS[1]), .B(HTRANS[0]), .C(HADDR[0]), .Y(n148) );
  NOR2X1 U242 ( .A(n149), .B(n150), .Y(n137) );
  NAND3X1 U243 ( .A(HADDR[11]), .B(HADDR[10]), .C(HADDR[12]), .Y(n150) );
  NAND3X1 U244 ( .A(HADDR[7]), .B(HADDR[6]), .C(HADDR[8]), .Y(n149) );
  AOI21X1 U247 ( .A(n153), .B(HTRANS[0]), .C(split), .Y(n152) );
  NOR2X1 U248 ( .A(HTRANS[1]), .B(HSEL), .Y(n153) );
  NOR2X1 U249 ( .A(n54), .B(n40), .Y(ADDR_RD[8]) );
  NOR2X1 U250 ( .A(n55), .B(n40), .Y(ADDR_RD[7]) );
  NOR2X1 U251 ( .A(n56), .B(n40), .Y(ADDR_RD[6]) );
  NOR2X1 U252 ( .A(n57), .B(n40), .Y(ADDR_RD[5]) );
  NOR2X1 U253 ( .A(n58), .B(n40), .Y(ADDR_RD[4]) );
  NOR2X1 U254 ( .A(n59), .B(n40), .Y(ADDR_RD[3]) );
  NOR2X1 U255 ( .A(n60), .B(n40), .Y(ADDR_RD[2]) );
  NOR2X1 U256 ( .A(n61), .B(n40), .Y(ADDR_RD[1]) );
  NOR2X1 U257 ( .A(n62), .B(n40), .Y(ADDR_RD[0]) );
  DFFSR \waitstate_pre_reg[1]  ( .D(N57), .CLK(clk), .R(n52), .S(1'b1), .Q(
        waitstate_pre[1]) );
  DFFSR \waitstate_pre_reg[0]  ( .D(N56), .CLK(clk), .R(n52), .S(1'b1), .Q(
        waitstate_pre[0]) );
  DFFSR \HSPLIT_reg[15]  ( .D(n165), .CLK(clk), .R(n52), .S(1'b1), .Q(
        HSPLIT[15]) );
  DFFSR \HSPLIT_reg[14]  ( .D(n166), .CLK(clk), .R(n52), .S(1'b1), .Q(
        HSPLIT[14]) );
  DFFSR \HSPLIT_reg[13]  ( .D(n167), .CLK(clk), .R(n52), .S(1'b1), .Q(
        HSPLIT[13]) );
  DFFSR \HSPLIT_reg[10]  ( .D(n170), .CLK(clk), .R(n52), .S(1'b1), .Q(
        HSPLIT[10]) );
  DFFSR \HSPLIT_reg[9]  ( .D(n171), .CLK(clk), .R(n52), .S(1'b1), .Q(HSPLIT[9]) );
  DFFSR \HSPLIT_reg[6]  ( .D(n174), .CLK(clk), .R(n52), .S(1'b1), .Q(HSPLIT[6]) );
  DFFSR \HSPLIT_reg[5]  ( .D(n175), .CLK(clk), .R(n52), .S(1'b1), .Q(HSPLIT[5]) );
  DFFSR \HSPLIT_reg[2]  ( .D(n178), .CLK(clk), .R(n52), .S(1'b1), .Q(HSPLIT[2]) );
  DFFSR \HSPLIT_reg[1]  ( .D(n179), .CLK(clk), .R(n52), .S(1'b1), .Q(HSPLIT[1]) );
  DFFSR \HRESP_reg[0]  ( .D(N34), .CLK(clk), .R(n52), .S(1'b1), .Q(HRESP[0])
         );
  DFFSR \HSPLIT_reg[12]  ( .D(n168), .CLK(clk), .R(n52), .S(1'b1), .Q(
        HSPLIT[12]) );
  DFFSR \HSPLIT_reg[11]  ( .D(n169), .CLK(clk), .R(n52), .S(1'b1), .Q(
        HSPLIT[11]) );
  DFFSR \HSPLIT_reg[8]  ( .D(n172), .CLK(clk), .R(n52), .S(1'b1), .Q(HSPLIT[8]) );
  DFFSR \HSPLIT_reg[7]  ( .D(n173), .CLK(clk), .R(n52), .S(1'b1), .Q(HSPLIT[7]) );
  DFFSR \HSPLIT_reg[4]  ( .D(n176), .CLK(clk), .R(n52), .S(1'b1), .Q(HSPLIT[4]) );
  DFFSR \HSPLIT_reg[3]  ( .D(n177), .CLK(clk), .R(n52), .S(1'b1), .Q(HSPLIT[3]) );
  DFFSR \HSPLIT_reg[0]  ( .D(n180), .CLK(clk), .R(n52), .S(1'b1), .Q(HSPLIT[0]) );
  DFFSR \HRESP_reg[1]  ( .D(n47), .CLK(clk), .R(n52), .S(1'b1), .Q(HRESP[1])
         );
  DFFSR \waitstate_reg[1]  ( .D(N36), .CLK(clk), .R(n52), .S(1'b1), .Q(
        waitstate[1]) );
  DFFSR split_reg ( .D(n181), .CLK(clk), .R(n52), .S(1'b1), .Q(split) );
  DFFSR \waitstate_reg[0]  ( .D(N35), .CLK(clk), .R(n52), .S(1'b1), .Q(
        waitstate[0]) );
  DFFSR \waitstate_reg[2]  ( .D(N37), .CLK(clk), .R(n52), .S(1'b1), .Q(
        waitstate[2]) );
  DFFSR data_phase_reg ( .D(n164), .CLK(clk), .R(n52), .S(1'b1), .Q(data_phase) );
  DFFSR WR_pre_d_reg ( .D(n154), .CLK(clk), .R(n52), .S(1'b1), .Q(WR_pre_d) );
  DFFSR \ADDR_WR_reg[8]  ( .D(n163), .CLK(clk), .R(n52), .S(1'b1), .Q(
        ADDR_WR[8]) );
  DFFSR \ADDR_WR_reg[7]  ( .D(n162), .CLK(clk), .R(n52), .S(1'b1), .Q(
        ADDR_WR[7]) );
  DFFSR \ADDR_WR_reg[6]  ( .D(n161), .CLK(clk), .R(n52), .S(1'b1), .Q(
        ADDR_WR[6]) );
  DFFSR \ADDR_WR_reg[5]  ( .D(n160), .CLK(clk), .R(n52), .S(1'b1), .Q(
        ADDR_WR[5]) );
  DFFSR \ADDR_WR_reg[4]  ( .D(n159), .CLK(clk), .R(n52), .S(1'b1), .Q(
        ADDR_WR[4]) );
  DFFSR \ADDR_WR_reg[3]  ( .D(n158), .CLK(clk), .R(n52), .S(1'b1), .Q(
        ADDR_WR[3]) );
  DFFSR \ADDR_WR_reg[2]  ( .D(n157), .CLK(clk), .R(n52), .S(1'b1), .Q(
        ADDR_WR[2]) );
  DFFSR \ADDR_WR_reg[1]  ( .D(n156), .CLK(clk), .R(n52), .S(1'b1), .Q(
        ADDR_WR[1]) );
  DFFSR \ADDR_WR_reg[0]  ( .D(n155), .CLK(clk), .R(n52), .S(1'b1), .Q(
        ADDR_WR[0]) );
  AND2X2 U3 ( .A(HTRANS[1]), .B(n64), .Y(RD) );
  AND2X2 U4 ( .A(n152), .B(STALL), .Y(n2) );
  XNOR2X1 U5 ( .A(waitstate_pre[0]), .B(waitstate[0]), .Y(n3) );
  INVX4 U6 ( .A(reset), .Y(n52) );
  INVX2 U115 ( .A(n46), .Y(HREADY) );
  INVX2 U116 ( .A(n39), .Y(n44) );
  INVX2 U117 ( .A(n2), .Y(n46) );
  BUFX2 U118 ( .A(n81), .Y(n41) );
  BUFX2 U119 ( .A(n81), .Y(n42) );
  OR2X2 U120 ( .A(n50), .B(n46), .Y(n39) );
  INVX2 U121 ( .A(RD), .Y(n40) );
  INVX2 U122 ( .A(n41), .Y(n47) );
  INVX2 U123 ( .A(waitstate[1]), .Y(n48) );
  INVX2 U124 ( .A(waitstate[2]), .Y(n49) );
  INVX2 U125 ( .A(data_phase), .Y(n50) );
  INVX2 U126 ( .A(WR_pre_d), .Y(n51) );
  INVX2 U127 ( .A(n104), .Y(n53) );
  INVX2 U128 ( .A(HADDR[8]), .Y(n54) );
  INVX2 U129 ( .A(HADDR[7]), .Y(n55) );
  INVX2 U130 ( .A(HADDR[6]), .Y(n56) );
  INVX2 U131 ( .A(HADDR[5]), .Y(n57) );
  INVX2 U132 ( .A(HADDR[4]), .Y(n58) );
  INVX2 U133 ( .A(HADDR[3]), .Y(n59) );
  INVX2 U134 ( .A(HADDR[2]), .Y(n60) );
  INVX2 U135 ( .A(HADDR[1]), .Y(n61) );
  INVX2 U136 ( .A(HADDR[0]), .Y(n62) );
  INVX2 U215 ( .A(n148), .Y(n63) );
  INVX2 U218 ( .A(HWRITE), .Y(n64) );
  INVX2 U219 ( .A(RANDSPLIT[2]), .Y(n65) );
  INVX2 U245 ( .A(HMASTER[2]), .Y(n66) );
  INVX2 U246 ( .A(HMASTER[1]), .Y(n67) );
  INVX2 U258 ( .A(HMASTER[0]), .Y(n70) );
endmodule


module ahb_slave_mem ( clk, reset, WR, RD, ADDR_WR, ADDR_RD, DIN, DOUT );
  input [8:0] ADDR_WR;
  input [8:0] ADDR_RD;
  input [31:0] DIN;
  output [31:0] DOUT;
  input clk, reset, WR, RD;
  wire   N10, N11, N12, N13, N14, N15, \Mem[63][31] , \Mem[63][30] ,
         \Mem[63][29] , \Mem[63][28] , \Mem[63][27] , \Mem[63][26] ,
         \Mem[63][25] , \Mem[63][24] , \Mem[63][23] , \Mem[63][22] ,
         \Mem[63][21] , \Mem[63][20] , \Mem[63][19] , \Mem[63][18] ,
         \Mem[63][17] , \Mem[63][16] , \Mem[63][15] , \Mem[63][14] ,
         \Mem[63][13] , \Mem[63][12] , \Mem[63][11] , \Mem[63][10] ,
         \Mem[63][9] , \Mem[63][8] , \Mem[63][7] , \Mem[63][6] , \Mem[63][5] ,
         \Mem[63][4] , \Mem[63][3] , \Mem[63][2] , \Mem[63][1] , \Mem[63][0] ,
         \Mem[62][31] , \Mem[62][30] , \Mem[62][29] , \Mem[62][28] ,
         \Mem[62][27] , \Mem[62][26] , \Mem[62][25] , \Mem[62][24] ,
         \Mem[62][23] , \Mem[62][22] , \Mem[62][21] , \Mem[62][20] ,
         \Mem[62][19] , \Mem[62][18] , \Mem[62][17] , \Mem[62][16] ,
         \Mem[62][15] , \Mem[62][14] , \Mem[62][13] , \Mem[62][12] ,
         \Mem[62][11] , \Mem[62][10] , \Mem[62][9] , \Mem[62][8] ,
         \Mem[62][7] , \Mem[62][6] , \Mem[62][5] , \Mem[62][4] , \Mem[62][3] ,
         \Mem[62][2] , \Mem[62][1] , \Mem[62][0] , \Mem[61][31] ,
         \Mem[61][30] , \Mem[61][29] , \Mem[61][28] , \Mem[61][27] ,
         \Mem[61][26] , \Mem[61][25] , \Mem[61][24] , \Mem[61][23] ,
         \Mem[61][22] , \Mem[61][21] , \Mem[61][20] , \Mem[61][19] ,
         \Mem[61][18] , \Mem[61][17] , \Mem[61][16] , \Mem[61][15] ,
         \Mem[61][14] , \Mem[61][13] , \Mem[61][12] , \Mem[61][11] ,
         \Mem[61][10] , \Mem[61][9] , \Mem[61][8] , \Mem[61][7] , \Mem[61][6] ,
         \Mem[61][5] , \Mem[61][4] , \Mem[61][3] , \Mem[61][2] , \Mem[61][1] ,
         \Mem[61][0] , \Mem[60][31] , \Mem[60][30] , \Mem[60][29] ,
         \Mem[60][28] , \Mem[60][27] , \Mem[60][26] , \Mem[60][25] ,
         \Mem[60][24] , \Mem[60][23] , \Mem[60][22] , \Mem[60][21] ,
         \Mem[60][20] , \Mem[60][19] , \Mem[60][18] , \Mem[60][17] ,
         \Mem[60][16] , \Mem[60][15] , \Mem[60][14] , \Mem[60][13] ,
         \Mem[60][12] , \Mem[60][11] , \Mem[60][10] , \Mem[60][9] ,
         \Mem[60][8] , \Mem[60][7] , \Mem[60][6] , \Mem[60][5] , \Mem[60][4] ,
         \Mem[60][3] , \Mem[60][2] , \Mem[60][1] , \Mem[60][0] , \Mem[59][31] ,
         \Mem[59][30] , \Mem[59][29] , \Mem[59][28] , \Mem[59][27] ,
         \Mem[59][26] , \Mem[59][25] , \Mem[59][24] , \Mem[59][23] ,
         \Mem[59][22] , \Mem[59][21] , \Mem[59][20] , \Mem[59][19] ,
         \Mem[59][18] , \Mem[59][17] , \Mem[59][16] , \Mem[59][15] ,
         \Mem[59][14] , \Mem[59][13] , \Mem[59][12] , \Mem[59][11] ,
         \Mem[59][10] , \Mem[59][9] , \Mem[59][8] , \Mem[59][7] , \Mem[59][6] ,
         \Mem[59][5] , \Mem[59][4] , \Mem[59][3] , \Mem[59][2] , \Mem[59][1] ,
         \Mem[59][0] , \Mem[58][31] , \Mem[58][30] , \Mem[58][29] ,
         \Mem[58][28] , \Mem[58][27] , \Mem[58][26] , \Mem[58][25] ,
         \Mem[58][24] , \Mem[58][23] , \Mem[58][22] , \Mem[58][21] ,
         \Mem[58][20] , \Mem[58][19] , \Mem[58][18] , \Mem[58][17] ,
         \Mem[58][16] , \Mem[58][15] , \Mem[58][14] , \Mem[58][13] ,
         \Mem[58][12] , \Mem[58][11] , \Mem[58][10] , \Mem[58][9] ,
         \Mem[58][8] , \Mem[58][7] , \Mem[58][6] , \Mem[58][5] , \Mem[58][4] ,
         \Mem[58][3] , \Mem[58][2] , \Mem[58][1] , \Mem[58][0] , \Mem[57][31] ,
         \Mem[57][30] , \Mem[57][29] , \Mem[57][28] , \Mem[57][27] ,
         \Mem[57][26] , \Mem[57][25] , \Mem[57][24] , \Mem[57][23] ,
         \Mem[57][22] , \Mem[57][21] , \Mem[57][20] , \Mem[57][19] ,
         \Mem[57][18] , \Mem[57][17] , \Mem[57][16] , \Mem[57][15] ,
         \Mem[57][14] , \Mem[57][13] , \Mem[57][12] , \Mem[57][11] ,
         \Mem[57][10] , \Mem[57][9] , \Mem[57][8] , \Mem[57][7] , \Mem[57][6] ,
         \Mem[57][5] , \Mem[57][4] , \Mem[57][3] , \Mem[57][2] , \Mem[57][1] ,
         \Mem[57][0] , \Mem[56][31] , \Mem[56][30] , \Mem[56][29] ,
         \Mem[56][28] , \Mem[56][27] , \Mem[56][26] , \Mem[56][25] ,
         \Mem[56][24] , \Mem[56][23] , \Mem[56][22] , \Mem[56][21] ,
         \Mem[56][20] , \Mem[56][19] , \Mem[56][18] , \Mem[56][17] ,
         \Mem[56][16] , \Mem[56][15] , \Mem[56][14] , \Mem[56][13] ,
         \Mem[56][12] , \Mem[56][11] , \Mem[56][10] , \Mem[56][9] ,
         \Mem[56][8] , \Mem[56][7] , \Mem[56][6] , \Mem[56][5] , \Mem[56][4] ,
         \Mem[56][3] , \Mem[56][2] , \Mem[56][1] , \Mem[56][0] , \Mem[55][31] ,
         \Mem[55][30] , \Mem[55][29] , \Mem[55][28] , \Mem[55][27] ,
         \Mem[55][26] , \Mem[55][25] , \Mem[55][24] , \Mem[55][23] ,
         \Mem[55][22] , \Mem[55][21] , \Mem[55][20] , \Mem[55][19] ,
         \Mem[55][18] , \Mem[55][17] , \Mem[55][16] , \Mem[55][15] ,
         \Mem[55][14] , \Mem[55][13] , \Mem[55][12] , \Mem[55][11] ,
         \Mem[55][10] , \Mem[55][9] , \Mem[55][8] , \Mem[55][7] , \Mem[55][6] ,
         \Mem[55][5] , \Mem[55][4] , \Mem[55][3] , \Mem[55][2] , \Mem[55][1] ,
         \Mem[55][0] , \Mem[54][31] , \Mem[54][30] , \Mem[54][29] ,
         \Mem[54][28] , \Mem[54][27] , \Mem[54][26] , \Mem[54][25] ,
         \Mem[54][24] , \Mem[54][23] , \Mem[54][22] , \Mem[54][21] ,
         \Mem[54][20] , \Mem[54][19] , \Mem[54][18] , \Mem[54][17] ,
         \Mem[54][16] , \Mem[54][15] , \Mem[54][14] , \Mem[54][13] ,
         \Mem[54][12] , \Mem[54][11] , \Mem[54][10] , \Mem[54][9] ,
         \Mem[54][8] , \Mem[54][7] , \Mem[54][6] , \Mem[54][5] , \Mem[54][4] ,
         \Mem[54][3] , \Mem[54][2] , \Mem[54][1] , \Mem[54][0] , \Mem[53][31] ,
         \Mem[53][30] , \Mem[53][29] , \Mem[53][28] , \Mem[53][27] ,
         \Mem[53][26] , \Mem[53][25] , \Mem[53][24] , \Mem[53][23] ,
         \Mem[53][22] , \Mem[53][21] , \Mem[53][20] , \Mem[53][19] ,
         \Mem[53][18] , \Mem[53][17] , \Mem[53][16] , \Mem[53][15] ,
         \Mem[53][14] , \Mem[53][13] , \Mem[53][12] , \Mem[53][11] ,
         \Mem[53][10] , \Mem[53][9] , \Mem[53][8] , \Mem[53][7] , \Mem[53][6] ,
         \Mem[53][5] , \Mem[53][4] , \Mem[53][3] , \Mem[53][2] , \Mem[53][1] ,
         \Mem[53][0] , \Mem[52][31] , \Mem[52][30] , \Mem[52][29] ,
         \Mem[52][28] , \Mem[52][27] , \Mem[52][26] , \Mem[52][25] ,
         \Mem[52][24] , \Mem[52][23] , \Mem[52][22] , \Mem[52][21] ,
         \Mem[52][20] , \Mem[52][19] , \Mem[52][18] , \Mem[52][17] ,
         \Mem[52][16] , \Mem[52][15] , \Mem[52][14] , \Mem[52][13] ,
         \Mem[52][12] , \Mem[52][11] , \Mem[52][10] , \Mem[52][9] ,
         \Mem[52][8] , \Mem[52][7] , \Mem[52][6] , \Mem[52][5] , \Mem[52][4] ,
         \Mem[52][3] , \Mem[52][2] , \Mem[52][1] , \Mem[52][0] , \Mem[51][31] ,
         \Mem[51][30] , \Mem[51][29] , \Mem[51][28] , \Mem[51][27] ,
         \Mem[51][26] , \Mem[51][25] , \Mem[51][24] , \Mem[51][23] ,
         \Mem[51][22] , \Mem[51][21] , \Mem[51][20] , \Mem[51][19] ,
         \Mem[51][18] , \Mem[51][17] , \Mem[51][16] , \Mem[51][15] ,
         \Mem[51][14] , \Mem[51][13] , \Mem[51][12] , \Mem[51][11] ,
         \Mem[51][10] , \Mem[51][9] , \Mem[51][8] , \Mem[51][7] , \Mem[51][6] ,
         \Mem[51][5] , \Mem[51][4] , \Mem[51][3] , \Mem[51][2] , \Mem[51][1] ,
         \Mem[51][0] , \Mem[50][31] , \Mem[50][30] , \Mem[50][29] ,
         \Mem[50][28] , \Mem[50][27] , \Mem[50][26] , \Mem[50][25] ,
         \Mem[50][24] , \Mem[50][23] , \Mem[50][22] , \Mem[50][21] ,
         \Mem[50][20] , \Mem[50][19] , \Mem[50][18] , \Mem[50][17] ,
         \Mem[50][16] , \Mem[50][15] , \Mem[50][14] , \Mem[50][13] ,
         \Mem[50][12] , \Mem[50][11] , \Mem[50][10] , \Mem[50][9] ,
         \Mem[50][8] , \Mem[50][7] , \Mem[50][6] , \Mem[50][5] , \Mem[50][4] ,
         \Mem[50][3] , \Mem[50][2] , \Mem[50][1] , \Mem[50][0] , \Mem[49][31] ,
         \Mem[49][30] , \Mem[49][29] , \Mem[49][28] , \Mem[49][27] ,
         \Mem[49][26] , \Mem[49][25] , \Mem[49][24] , \Mem[49][23] ,
         \Mem[49][22] , \Mem[49][21] , \Mem[49][20] , \Mem[49][19] ,
         \Mem[49][18] , \Mem[49][17] , \Mem[49][16] , \Mem[49][15] ,
         \Mem[49][14] , \Mem[49][13] , \Mem[49][12] , \Mem[49][11] ,
         \Mem[49][10] , \Mem[49][9] , \Mem[49][8] , \Mem[49][7] , \Mem[49][6] ,
         \Mem[49][5] , \Mem[49][4] , \Mem[49][3] , \Mem[49][2] , \Mem[49][1] ,
         \Mem[49][0] , \Mem[48][31] , \Mem[48][30] , \Mem[48][29] ,
         \Mem[48][28] , \Mem[48][27] , \Mem[48][26] , \Mem[48][25] ,
         \Mem[48][24] , \Mem[48][23] , \Mem[48][22] , \Mem[48][21] ,
         \Mem[48][20] , \Mem[48][19] , \Mem[48][18] , \Mem[48][17] ,
         \Mem[48][16] , \Mem[48][15] , \Mem[48][14] , \Mem[48][13] ,
         \Mem[48][12] , \Mem[48][11] , \Mem[48][10] , \Mem[48][9] ,
         \Mem[48][8] , \Mem[48][7] , \Mem[48][6] , \Mem[48][5] , \Mem[48][4] ,
         \Mem[48][3] , \Mem[48][2] , \Mem[48][1] , \Mem[48][0] , \Mem[47][31] ,
         \Mem[47][30] , \Mem[47][29] , \Mem[47][28] , \Mem[47][27] ,
         \Mem[47][26] , \Mem[47][25] , \Mem[47][24] , \Mem[47][23] ,
         \Mem[47][22] , \Mem[47][21] , \Mem[47][20] , \Mem[47][19] ,
         \Mem[47][18] , \Mem[47][17] , \Mem[47][16] , \Mem[47][15] ,
         \Mem[47][14] , \Mem[47][13] , \Mem[47][12] , \Mem[47][11] ,
         \Mem[47][10] , \Mem[47][9] , \Mem[47][8] , \Mem[47][7] , \Mem[47][6] ,
         \Mem[47][5] , \Mem[47][4] , \Mem[47][3] , \Mem[47][2] , \Mem[47][1] ,
         \Mem[47][0] , \Mem[46][31] , \Mem[46][30] , \Mem[46][29] ,
         \Mem[46][28] , \Mem[46][27] , \Mem[46][26] , \Mem[46][25] ,
         \Mem[46][24] , \Mem[46][23] , \Mem[46][22] , \Mem[46][21] ,
         \Mem[46][20] , \Mem[46][19] , \Mem[46][18] , \Mem[46][17] ,
         \Mem[46][16] , \Mem[46][15] , \Mem[46][14] , \Mem[46][13] ,
         \Mem[46][12] , \Mem[46][11] , \Mem[46][10] , \Mem[46][9] ,
         \Mem[46][8] , \Mem[46][7] , \Mem[46][6] , \Mem[46][5] , \Mem[46][4] ,
         \Mem[46][3] , \Mem[46][2] , \Mem[46][1] , \Mem[46][0] , \Mem[45][31] ,
         \Mem[45][30] , \Mem[45][29] , \Mem[45][28] , \Mem[45][27] ,
         \Mem[45][26] , \Mem[45][25] , \Mem[45][24] , \Mem[45][23] ,
         \Mem[45][22] , \Mem[45][21] , \Mem[45][20] , \Mem[45][19] ,
         \Mem[45][18] , \Mem[45][17] , \Mem[45][16] , \Mem[45][15] ,
         \Mem[45][14] , \Mem[45][13] , \Mem[45][12] , \Mem[45][11] ,
         \Mem[45][10] , \Mem[45][9] , \Mem[45][8] , \Mem[45][7] , \Mem[45][6] ,
         \Mem[45][5] , \Mem[45][4] , \Mem[45][3] , \Mem[45][2] , \Mem[45][1] ,
         \Mem[45][0] , \Mem[44][31] , \Mem[44][30] , \Mem[44][29] ,
         \Mem[44][28] , \Mem[44][27] , \Mem[44][26] , \Mem[44][25] ,
         \Mem[44][24] , \Mem[44][23] , \Mem[44][22] , \Mem[44][21] ,
         \Mem[44][20] , \Mem[44][19] , \Mem[44][18] , \Mem[44][17] ,
         \Mem[44][16] , \Mem[44][15] , \Mem[44][14] , \Mem[44][13] ,
         \Mem[44][12] , \Mem[44][11] , \Mem[44][10] , \Mem[44][9] ,
         \Mem[44][8] , \Mem[44][7] , \Mem[44][6] , \Mem[44][5] , \Mem[44][4] ,
         \Mem[44][3] , \Mem[44][2] , \Mem[44][1] , \Mem[44][0] , \Mem[43][31] ,
         \Mem[43][30] , \Mem[43][29] , \Mem[43][28] , \Mem[43][27] ,
         \Mem[43][26] , \Mem[43][25] , \Mem[43][24] , \Mem[43][23] ,
         \Mem[43][22] , \Mem[43][21] , \Mem[43][20] , \Mem[43][19] ,
         \Mem[43][18] , \Mem[43][17] , \Mem[43][16] , \Mem[43][15] ,
         \Mem[43][14] , \Mem[43][13] , \Mem[43][12] , \Mem[43][11] ,
         \Mem[43][10] , \Mem[43][9] , \Mem[43][8] , \Mem[43][7] , \Mem[43][6] ,
         \Mem[43][5] , \Mem[43][4] , \Mem[43][3] , \Mem[43][2] , \Mem[43][1] ,
         \Mem[43][0] , \Mem[42][31] , \Mem[42][30] , \Mem[42][29] ,
         \Mem[42][28] , \Mem[42][27] , \Mem[42][26] , \Mem[42][25] ,
         \Mem[42][24] , \Mem[42][23] , \Mem[42][22] , \Mem[42][21] ,
         \Mem[42][20] , \Mem[42][19] , \Mem[42][18] , \Mem[42][17] ,
         \Mem[42][16] , \Mem[42][15] , \Mem[42][14] , \Mem[42][13] ,
         \Mem[42][12] , \Mem[42][11] , \Mem[42][10] , \Mem[42][9] ,
         \Mem[42][8] , \Mem[42][7] , \Mem[42][6] , \Mem[42][5] , \Mem[42][4] ,
         \Mem[42][3] , \Mem[42][2] , \Mem[42][1] , \Mem[42][0] , \Mem[41][31] ,
         \Mem[41][30] , \Mem[41][29] , \Mem[41][28] , \Mem[41][27] ,
         \Mem[41][26] , \Mem[41][25] , \Mem[41][24] , \Mem[41][23] ,
         \Mem[41][22] , \Mem[41][21] , \Mem[41][20] , \Mem[41][19] ,
         \Mem[41][18] , \Mem[41][17] , \Mem[41][16] , \Mem[41][15] ,
         \Mem[41][14] , \Mem[41][13] , \Mem[41][12] , \Mem[41][11] ,
         \Mem[41][10] , \Mem[41][9] , \Mem[41][8] , \Mem[41][7] , \Mem[41][6] ,
         \Mem[41][5] , \Mem[41][4] , \Mem[41][3] , \Mem[41][2] , \Mem[41][1] ,
         \Mem[41][0] , \Mem[40][31] , \Mem[40][30] , \Mem[40][29] ,
         \Mem[40][28] , \Mem[40][27] , \Mem[40][26] , \Mem[40][25] ,
         \Mem[40][24] , \Mem[40][23] , \Mem[40][22] , \Mem[40][21] ,
         \Mem[40][20] , \Mem[40][19] , \Mem[40][18] , \Mem[40][17] ,
         \Mem[40][16] , \Mem[40][15] , \Mem[40][14] , \Mem[40][13] ,
         \Mem[40][12] , \Mem[40][11] , \Mem[40][10] , \Mem[40][9] ,
         \Mem[40][8] , \Mem[40][7] , \Mem[40][6] , \Mem[40][5] , \Mem[40][4] ,
         \Mem[40][3] , \Mem[40][2] , \Mem[40][1] , \Mem[40][0] , \Mem[39][31] ,
         \Mem[39][30] , \Mem[39][29] , \Mem[39][28] , \Mem[39][27] ,
         \Mem[39][26] , \Mem[39][25] , \Mem[39][24] , \Mem[39][23] ,
         \Mem[39][22] , \Mem[39][21] , \Mem[39][20] , \Mem[39][19] ,
         \Mem[39][18] , \Mem[39][17] , \Mem[39][16] , \Mem[39][15] ,
         \Mem[39][14] , \Mem[39][13] , \Mem[39][12] , \Mem[39][11] ,
         \Mem[39][10] , \Mem[39][9] , \Mem[39][8] , \Mem[39][7] , \Mem[39][6] ,
         \Mem[39][5] , \Mem[39][4] , \Mem[39][3] , \Mem[39][2] , \Mem[39][1] ,
         \Mem[39][0] , \Mem[38][31] , \Mem[38][30] , \Mem[38][29] ,
         \Mem[38][28] , \Mem[38][27] , \Mem[38][26] , \Mem[38][25] ,
         \Mem[38][24] , \Mem[38][23] , \Mem[38][22] , \Mem[38][21] ,
         \Mem[38][20] , \Mem[38][19] , \Mem[38][18] , \Mem[38][17] ,
         \Mem[38][16] , \Mem[38][15] , \Mem[38][14] , \Mem[38][13] ,
         \Mem[38][12] , \Mem[38][11] , \Mem[38][10] , \Mem[38][9] ,
         \Mem[38][8] , \Mem[38][7] , \Mem[38][6] , \Mem[38][5] , \Mem[38][4] ,
         \Mem[38][3] , \Mem[38][2] , \Mem[38][1] , \Mem[38][0] , \Mem[37][31] ,
         \Mem[37][30] , \Mem[37][29] , \Mem[37][28] , \Mem[37][27] ,
         \Mem[37][26] , \Mem[37][25] , \Mem[37][24] , \Mem[37][23] ,
         \Mem[37][22] , \Mem[37][21] , \Mem[37][20] , \Mem[37][19] ,
         \Mem[37][18] , \Mem[37][17] , \Mem[37][16] , \Mem[37][15] ,
         \Mem[37][14] , \Mem[37][13] , \Mem[37][12] , \Mem[37][11] ,
         \Mem[37][10] , \Mem[37][9] , \Mem[37][8] , \Mem[37][7] , \Mem[37][6] ,
         \Mem[37][5] , \Mem[37][4] , \Mem[37][3] , \Mem[37][2] , \Mem[37][1] ,
         \Mem[37][0] , \Mem[36][31] , \Mem[36][30] , \Mem[36][29] ,
         \Mem[36][28] , \Mem[36][27] , \Mem[36][26] , \Mem[36][25] ,
         \Mem[36][24] , \Mem[36][23] , \Mem[36][22] , \Mem[36][21] ,
         \Mem[36][20] , \Mem[36][19] , \Mem[36][18] , \Mem[36][17] ,
         \Mem[36][16] , \Mem[36][15] , \Mem[36][14] , \Mem[36][13] ,
         \Mem[36][12] , \Mem[36][11] , \Mem[36][10] , \Mem[36][9] ,
         \Mem[36][8] , \Mem[36][7] , \Mem[36][6] , \Mem[36][5] , \Mem[36][4] ,
         \Mem[36][3] , \Mem[36][2] , \Mem[36][1] , \Mem[36][0] , \Mem[35][31] ,
         \Mem[35][30] , \Mem[35][29] , \Mem[35][28] , \Mem[35][27] ,
         \Mem[35][26] , \Mem[35][25] , \Mem[35][24] , \Mem[35][23] ,
         \Mem[35][22] , \Mem[35][21] , \Mem[35][20] , \Mem[35][19] ,
         \Mem[35][18] , \Mem[35][17] , \Mem[35][16] , \Mem[35][15] ,
         \Mem[35][14] , \Mem[35][13] , \Mem[35][12] , \Mem[35][11] ,
         \Mem[35][10] , \Mem[35][9] , \Mem[35][8] , \Mem[35][7] , \Mem[35][6] ,
         \Mem[35][5] , \Mem[35][4] , \Mem[35][3] , \Mem[35][2] , \Mem[35][1] ,
         \Mem[35][0] , \Mem[34][31] , \Mem[34][30] , \Mem[34][29] ,
         \Mem[34][28] , \Mem[34][27] , \Mem[34][26] , \Mem[34][25] ,
         \Mem[34][24] , \Mem[34][23] , \Mem[34][22] , \Mem[34][21] ,
         \Mem[34][20] , \Mem[34][19] , \Mem[34][18] , \Mem[34][17] ,
         \Mem[34][16] , \Mem[34][15] , \Mem[34][14] , \Mem[34][13] ,
         \Mem[34][12] , \Mem[34][11] , \Mem[34][10] , \Mem[34][9] ,
         \Mem[34][8] , \Mem[34][7] , \Mem[34][6] , \Mem[34][5] , \Mem[34][4] ,
         \Mem[34][3] , \Mem[34][2] , \Mem[34][1] , \Mem[34][0] , \Mem[33][31] ,
         \Mem[33][30] , \Mem[33][29] , \Mem[33][28] , \Mem[33][27] ,
         \Mem[33][26] , \Mem[33][25] , \Mem[33][24] , \Mem[33][23] ,
         \Mem[33][22] , \Mem[33][21] , \Mem[33][20] , \Mem[33][19] ,
         \Mem[33][18] , \Mem[33][17] , \Mem[33][16] , \Mem[33][15] ,
         \Mem[33][14] , \Mem[33][13] , \Mem[33][12] , \Mem[33][11] ,
         \Mem[33][10] , \Mem[33][9] , \Mem[33][8] , \Mem[33][7] , \Mem[33][6] ,
         \Mem[33][5] , \Mem[33][4] , \Mem[33][3] , \Mem[33][2] , \Mem[33][1] ,
         \Mem[33][0] , \Mem[32][31] , \Mem[32][30] , \Mem[32][29] ,
         \Mem[32][28] , \Mem[32][27] , \Mem[32][26] , \Mem[32][25] ,
         \Mem[32][24] , \Mem[32][23] , \Mem[32][22] , \Mem[32][21] ,
         \Mem[32][20] , \Mem[32][19] , \Mem[32][18] , \Mem[32][17] ,
         \Mem[32][16] , \Mem[32][15] , \Mem[32][14] , \Mem[32][13] ,
         \Mem[32][12] , \Mem[32][11] , \Mem[32][10] , \Mem[32][9] ,
         \Mem[32][8] , \Mem[32][7] , \Mem[32][6] , \Mem[32][5] , \Mem[32][4] ,
         \Mem[32][3] , \Mem[32][2] , \Mem[32][1] , \Mem[32][0] , \Mem[31][31] ,
         \Mem[31][30] , \Mem[31][29] , \Mem[31][28] , \Mem[31][27] ,
         \Mem[31][26] , \Mem[31][25] , \Mem[31][24] , \Mem[31][23] ,
         \Mem[31][22] , \Mem[31][21] , \Mem[31][20] , \Mem[31][19] ,
         \Mem[31][18] , \Mem[31][17] , \Mem[31][16] , \Mem[31][15] ,
         \Mem[31][14] , \Mem[31][13] , \Mem[31][12] , \Mem[31][11] ,
         \Mem[31][10] , \Mem[31][9] , \Mem[31][8] , \Mem[31][7] , \Mem[31][6] ,
         \Mem[31][5] , \Mem[31][4] , \Mem[31][3] , \Mem[31][2] , \Mem[31][1] ,
         \Mem[31][0] , \Mem[30][31] , \Mem[30][30] , \Mem[30][29] ,
         \Mem[30][28] , \Mem[30][27] , \Mem[30][26] , \Mem[30][25] ,
         \Mem[30][24] , \Mem[30][23] , \Mem[30][22] , \Mem[30][21] ,
         \Mem[30][20] , \Mem[30][19] , \Mem[30][18] , \Mem[30][17] ,
         \Mem[30][16] , \Mem[30][15] , \Mem[30][14] , \Mem[30][13] ,
         \Mem[30][12] , \Mem[30][11] , \Mem[30][10] , \Mem[30][9] ,
         \Mem[30][8] , \Mem[30][7] , \Mem[30][6] , \Mem[30][5] , \Mem[30][4] ,
         \Mem[30][3] , \Mem[30][2] , \Mem[30][1] , \Mem[30][0] , \Mem[29][31] ,
         \Mem[29][30] , \Mem[29][29] , \Mem[29][28] , \Mem[29][27] ,
         \Mem[29][26] , \Mem[29][25] , \Mem[29][24] , \Mem[29][23] ,
         \Mem[29][22] , \Mem[29][21] , \Mem[29][20] , \Mem[29][19] ,
         \Mem[29][18] , \Mem[29][17] , \Mem[29][16] , \Mem[29][15] ,
         \Mem[29][14] , \Mem[29][13] , \Mem[29][12] , \Mem[29][11] ,
         \Mem[29][10] , \Mem[29][9] , \Mem[29][8] , \Mem[29][7] , \Mem[29][6] ,
         \Mem[29][5] , \Mem[29][4] , \Mem[29][3] , \Mem[29][2] , \Mem[29][1] ,
         \Mem[29][0] , \Mem[28][31] , \Mem[28][30] , \Mem[28][29] ,
         \Mem[28][28] , \Mem[28][27] , \Mem[28][26] , \Mem[28][25] ,
         \Mem[28][24] , \Mem[28][23] , \Mem[28][22] , \Mem[28][21] ,
         \Mem[28][20] , \Mem[28][19] , \Mem[28][18] , \Mem[28][17] ,
         \Mem[28][16] , \Mem[28][15] , \Mem[28][14] , \Mem[28][13] ,
         \Mem[28][12] , \Mem[28][11] , \Mem[28][10] , \Mem[28][9] ,
         \Mem[28][8] , \Mem[28][7] , \Mem[28][6] , \Mem[28][5] , \Mem[28][4] ,
         \Mem[28][3] , \Mem[28][2] , \Mem[28][1] , \Mem[28][0] , \Mem[27][31] ,
         \Mem[27][30] , \Mem[27][29] , \Mem[27][28] , \Mem[27][27] ,
         \Mem[27][26] , \Mem[27][25] , \Mem[27][24] , \Mem[27][23] ,
         \Mem[27][22] , \Mem[27][21] , \Mem[27][20] , \Mem[27][19] ,
         \Mem[27][18] , \Mem[27][17] , \Mem[27][16] , \Mem[27][15] ,
         \Mem[27][14] , \Mem[27][13] , \Mem[27][12] , \Mem[27][11] ,
         \Mem[27][10] , \Mem[27][9] , \Mem[27][8] , \Mem[27][7] , \Mem[27][6] ,
         \Mem[27][5] , \Mem[27][4] , \Mem[27][3] , \Mem[27][2] , \Mem[27][1] ,
         \Mem[27][0] , \Mem[26][31] , \Mem[26][30] , \Mem[26][29] ,
         \Mem[26][28] , \Mem[26][27] , \Mem[26][26] , \Mem[26][25] ,
         \Mem[26][24] , \Mem[26][23] , \Mem[26][22] , \Mem[26][21] ,
         \Mem[26][20] , \Mem[26][19] , \Mem[26][18] , \Mem[26][17] ,
         \Mem[26][16] , \Mem[26][15] , \Mem[26][14] , \Mem[26][13] ,
         \Mem[26][12] , \Mem[26][11] , \Mem[26][10] , \Mem[26][9] ,
         \Mem[26][8] , \Mem[26][7] , \Mem[26][6] , \Mem[26][5] , \Mem[26][4] ,
         \Mem[26][3] , \Mem[26][2] , \Mem[26][1] , \Mem[26][0] , \Mem[25][31] ,
         \Mem[25][30] , \Mem[25][29] , \Mem[25][28] , \Mem[25][27] ,
         \Mem[25][26] , \Mem[25][25] , \Mem[25][24] , \Mem[25][23] ,
         \Mem[25][22] , \Mem[25][21] , \Mem[25][20] , \Mem[25][19] ,
         \Mem[25][18] , \Mem[25][17] , \Mem[25][16] , \Mem[25][15] ,
         \Mem[25][14] , \Mem[25][13] , \Mem[25][12] , \Mem[25][11] ,
         \Mem[25][10] , \Mem[25][9] , \Mem[25][8] , \Mem[25][7] , \Mem[25][6] ,
         \Mem[25][5] , \Mem[25][4] , \Mem[25][3] , \Mem[25][2] , \Mem[25][1] ,
         \Mem[25][0] , \Mem[24][31] , \Mem[24][30] , \Mem[24][29] ,
         \Mem[24][28] , \Mem[24][27] , \Mem[24][26] , \Mem[24][25] ,
         \Mem[24][24] , \Mem[24][23] , \Mem[24][22] , \Mem[24][21] ,
         \Mem[24][20] , \Mem[24][19] , \Mem[24][18] , \Mem[24][17] ,
         \Mem[24][16] , \Mem[24][15] , \Mem[24][14] , \Mem[24][13] ,
         \Mem[24][12] , \Mem[24][11] , \Mem[24][10] , \Mem[24][9] ,
         \Mem[24][8] , \Mem[24][7] , \Mem[24][6] , \Mem[24][5] , \Mem[24][4] ,
         \Mem[24][3] , \Mem[24][2] , \Mem[24][1] , \Mem[24][0] , \Mem[23][31] ,
         \Mem[23][30] , \Mem[23][29] , \Mem[23][28] , \Mem[23][27] ,
         \Mem[23][26] , \Mem[23][25] , \Mem[23][24] , \Mem[23][23] ,
         \Mem[23][22] , \Mem[23][21] , \Mem[23][20] , \Mem[23][19] ,
         \Mem[23][18] , \Mem[23][17] , \Mem[23][16] , \Mem[23][15] ,
         \Mem[23][14] , \Mem[23][13] , \Mem[23][12] , \Mem[23][11] ,
         \Mem[23][10] , \Mem[23][9] , \Mem[23][8] , \Mem[23][7] , \Mem[23][6] ,
         \Mem[23][5] , \Mem[23][4] , \Mem[23][3] , \Mem[23][2] , \Mem[23][1] ,
         \Mem[23][0] , \Mem[22][31] , \Mem[22][30] , \Mem[22][29] ,
         \Mem[22][28] , \Mem[22][27] , \Mem[22][26] , \Mem[22][25] ,
         \Mem[22][24] , \Mem[22][23] , \Mem[22][22] , \Mem[22][21] ,
         \Mem[22][20] , \Mem[22][19] , \Mem[22][18] , \Mem[22][17] ,
         \Mem[22][16] , \Mem[22][15] , \Mem[22][14] , \Mem[22][13] ,
         \Mem[22][12] , \Mem[22][11] , \Mem[22][10] , \Mem[22][9] ,
         \Mem[22][8] , \Mem[22][7] , \Mem[22][6] , \Mem[22][5] , \Mem[22][4] ,
         \Mem[22][3] , \Mem[22][2] , \Mem[22][1] , \Mem[22][0] , \Mem[21][31] ,
         \Mem[21][30] , \Mem[21][29] , \Mem[21][28] , \Mem[21][27] ,
         \Mem[21][26] , \Mem[21][25] , \Mem[21][24] , \Mem[21][23] ,
         \Mem[21][22] , \Mem[21][21] , \Mem[21][20] , \Mem[21][19] ,
         \Mem[21][18] , \Mem[21][17] , \Mem[21][16] , \Mem[21][15] ,
         \Mem[21][14] , \Mem[21][13] , \Mem[21][12] , \Mem[21][11] ,
         \Mem[21][10] , \Mem[21][9] , \Mem[21][8] , \Mem[21][7] , \Mem[21][6] ,
         \Mem[21][5] , \Mem[21][4] , \Mem[21][3] , \Mem[21][2] , \Mem[21][1] ,
         \Mem[21][0] , \Mem[20][31] , \Mem[20][30] , \Mem[20][29] ,
         \Mem[20][28] , \Mem[20][27] , \Mem[20][26] , \Mem[20][25] ,
         \Mem[20][24] , \Mem[20][23] , \Mem[20][22] , \Mem[20][21] ,
         \Mem[20][20] , \Mem[20][19] , \Mem[20][18] , \Mem[20][17] ,
         \Mem[20][16] , \Mem[20][15] , \Mem[20][14] , \Mem[20][13] ,
         \Mem[20][12] , \Mem[20][11] , \Mem[20][10] , \Mem[20][9] ,
         \Mem[20][8] , \Mem[20][7] , \Mem[20][6] , \Mem[20][5] , \Mem[20][4] ,
         \Mem[20][3] , \Mem[20][2] , \Mem[20][1] , \Mem[20][0] , \Mem[19][31] ,
         \Mem[19][30] , \Mem[19][29] , \Mem[19][28] , \Mem[19][27] ,
         \Mem[19][26] , \Mem[19][25] , \Mem[19][24] , \Mem[19][23] ,
         \Mem[19][22] , \Mem[19][21] , \Mem[19][20] , \Mem[19][19] ,
         \Mem[19][18] , \Mem[19][17] , \Mem[19][16] , \Mem[19][15] ,
         \Mem[19][14] , \Mem[19][13] , \Mem[19][12] , \Mem[19][11] ,
         \Mem[19][10] , \Mem[19][9] , \Mem[19][8] , \Mem[19][7] , \Mem[19][6] ,
         \Mem[19][5] , \Mem[19][4] , \Mem[19][3] , \Mem[19][2] , \Mem[19][1] ,
         \Mem[19][0] , \Mem[18][31] , \Mem[18][30] , \Mem[18][29] ,
         \Mem[18][28] , \Mem[18][27] , \Mem[18][26] , \Mem[18][25] ,
         \Mem[18][24] , \Mem[18][23] , \Mem[18][22] , \Mem[18][21] ,
         \Mem[18][20] , \Mem[18][19] , \Mem[18][18] , \Mem[18][17] ,
         \Mem[18][16] , \Mem[18][15] , \Mem[18][14] , \Mem[18][13] ,
         \Mem[18][12] , \Mem[18][11] , \Mem[18][10] , \Mem[18][9] ,
         \Mem[18][8] , \Mem[18][7] , \Mem[18][6] , \Mem[18][5] , \Mem[18][4] ,
         \Mem[18][3] , \Mem[18][2] , \Mem[18][1] , \Mem[18][0] , \Mem[17][31] ,
         \Mem[17][30] , \Mem[17][29] , \Mem[17][28] , \Mem[17][27] ,
         \Mem[17][26] , \Mem[17][25] , \Mem[17][24] , \Mem[17][23] ,
         \Mem[17][22] , \Mem[17][21] , \Mem[17][20] , \Mem[17][19] ,
         \Mem[17][18] , \Mem[17][17] , \Mem[17][16] , \Mem[17][15] ,
         \Mem[17][14] , \Mem[17][13] , \Mem[17][12] , \Mem[17][11] ,
         \Mem[17][10] , \Mem[17][9] , \Mem[17][8] , \Mem[17][7] , \Mem[17][6] ,
         \Mem[17][5] , \Mem[17][4] , \Mem[17][3] , \Mem[17][2] , \Mem[17][1] ,
         \Mem[17][0] , \Mem[16][31] , \Mem[16][30] , \Mem[16][29] ,
         \Mem[16][28] , \Mem[16][27] , \Mem[16][26] , \Mem[16][25] ,
         \Mem[16][24] , \Mem[16][23] , \Mem[16][22] , \Mem[16][21] ,
         \Mem[16][20] , \Mem[16][19] , \Mem[16][18] , \Mem[16][17] ,
         \Mem[16][16] , \Mem[16][15] , \Mem[16][14] , \Mem[16][13] ,
         \Mem[16][12] , \Mem[16][11] , \Mem[16][10] , \Mem[16][9] ,
         \Mem[16][8] , \Mem[16][7] , \Mem[16][6] , \Mem[16][5] , \Mem[16][4] ,
         \Mem[16][3] , \Mem[16][2] , \Mem[16][1] , \Mem[16][0] , \Mem[15][31] ,
         \Mem[15][30] , \Mem[15][29] , \Mem[15][28] , \Mem[15][27] ,
         \Mem[15][26] , \Mem[15][25] , \Mem[15][24] , \Mem[15][23] ,
         \Mem[15][22] , \Mem[15][21] , \Mem[15][20] , \Mem[15][19] ,
         \Mem[15][18] , \Mem[15][17] , \Mem[15][16] , \Mem[15][15] ,
         \Mem[15][14] , \Mem[15][13] , \Mem[15][12] , \Mem[15][11] ,
         \Mem[15][10] , \Mem[15][9] , \Mem[15][8] , \Mem[15][7] , \Mem[15][6] ,
         \Mem[15][5] , \Mem[15][4] , \Mem[15][3] , \Mem[15][2] , \Mem[15][1] ,
         \Mem[15][0] , \Mem[14][31] , \Mem[14][30] , \Mem[14][29] ,
         \Mem[14][28] , \Mem[14][27] , \Mem[14][26] , \Mem[14][25] ,
         \Mem[14][24] , \Mem[14][23] , \Mem[14][22] , \Mem[14][21] ,
         \Mem[14][20] , \Mem[14][19] , \Mem[14][18] , \Mem[14][17] ,
         \Mem[14][16] , \Mem[14][15] , \Mem[14][14] , \Mem[14][13] ,
         \Mem[14][12] , \Mem[14][11] , \Mem[14][10] , \Mem[14][9] ,
         \Mem[14][8] , \Mem[14][7] , \Mem[14][6] , \Mem[14][5] , \Mem[14][4] ,
         \Mem[14][3] , \Mem[14][2] , \Mem[14][1] , \Mem[14][0] , \Mem[13][31] ,
         \Mem[13][30] , \Mem[13][29] , \Mem[13][28] , \Mem[13][27] ,
         \Mem[13][26] , \Mem[13][25] , \Mem[13][24] , \Mem[13][23] ,
         \Mem[13][22] , \Mem[13][21] , \Mem[13][20] , \Mem[13][19] ,
         \Mem[13][18] , \Mem[13][17] , \Mem[13][16] , \Mem[13][15] ,
         \Mem[13][14] , \Mem[13][13] , \Mem[13][12] , \Mem[13][11] ,
         \Mem[13][10] , \Mem[13][9] , \Mem[13][8] , \Mem[13][7] , \Mem[13][6] ,
         \Mem[13][5] , \Mem[13][4] , \Mem[13][3] , \Mem[13][2] , \Mem[13][1] ,
         \Mem[13][0] , \Mem[12][31] , \Mem[12][30] , \Mem[12][29] ,
         \Mem[12][28] , \Mem[12][27] , \Mem[12][26] , \Mem[12][25] ,
         \Mem[12][24] , \Mem[12][23] , \Mem[12][22] , \Mem[12][21] ,
         \Mem[12][20] , \Mem[12][19] , \Mem[12][18] , \Mem[12][17] ,
         \Mem[12][16] , \Mem[12][15] , \Mem[12][14] , \Mem[12][13] ,
         \Mem[12][12] , \Mem[12][11] , \Mem[12][10] , \Mem[12][9] ,
         \Mem[12][8] , \Mem[12][7] , \Mem[12][6] , \Mem[12][5] , \Mem[12][4] ,
         \Mem[12][3] , \Mem[12][2] , \Mem[12][1] , \Mem[12][0] , \Mem[11][31] ,
         \Mem[11][30] , \Mem[11][29] , \Mem[11][28] , \Mem[11][27] ,
         \Mem[11][26] , \Mem[11][25] , \Mem[11][24] , \Mem[11][23] ,
         \Mem[11][22] , \Mem[11][21] , \Mem[11][20] , \Mem[11][19] ,
         \Mem[11][18] , \Mem[11][17] , \Mem[11][16] , \Mem[11][15] ,
         \Mem[11][14] , \Mem[11][13] , \Mem[11][12] , \Mem[11][11] ,
         \Mem[11][10] , \Mem[11][9] , \Mem[11][8] , \Mem[11][7] , \Mem[11][6] ,
         \Mem[11][5] , \Mem[11][4] , \Mem[11][3] , \Mem[11][2] , \Mem[11][1] ,
         \Mem[11][0] , \Mem[10][31] , \Mem[10][30] , \Mem[10][29] ,
         \Mem[10][28] , \Mem[10][27] , \Mem[10][26] , \Mem[10][25] ,
         \Mem[10][24] , \Mem[10][23] , \Mem[10][22] , \Mem[10][21] ,
         \Mem[10][20] , \Mem[10][19] , \Mem[10][18] , \Mem[10][17] ,
         \Mem[10][16] , \Mem[10][15] , \Mem[10][14] , \Mem[10][13] ,
         \Mem[10][12] , \Mem[10][11] , \Mem[10][10] , \Mem[10][9] ,
         \Mem[10][8] , \Mem[10][7] , \Mem[10][6] , \Mem[10][5] , \Mem[10][4] ,
         \Mem[10][3] , \Mem[10][2] , \Mem[10][1] , \Mem[10][0] , \Mem[9][31] ,
         \Mem[9][30] , \Mem[9][29] , \Mem[9][28] , \Mem[9][27] , \Mem[9][26] ,
         \Mem[9][25] , \Mem[9][24] , \Mem[9][23] , \Mem[9][22] , \Mem[9][21] ,
         \Mem[9][20] , \Mem[9][19] , \Mem[9][18] , \Mem[9][17] , \Mem[9][16] ,
         \Mem[9][15] , \Mem[9][14] , \Mem[9][13] , \Mem[9][12] , \Mem[9][11] ,
         \Mem[9][10] , \Mem[9][9] , \Mem[9][8] , \Mem[9][7] , \Mem[9][6] ,
         \Mem[9][5] , \Mem[9][4] , \Mem[9][3] , \Mem[9][2] , \Mem[9][1] ,
         \Mem[9][0] , \Mem[8][31] , \Mem[8][30] , \Mem[8][29] , \Mem[8][28] ,
         \Mem[8][27] , \Mem[8][26] , \Mem[8][25] , \Mem[8][24] , \Mem[8][23] ,
         \Mem[8][22] , \Mem[8][21] , \Mem[8][20] , \Mem[8][19] , \Mem[8][18] ,
         \Mem[8][17] , \Mem[8][16] , \Mem[8][15] , \Mem[8][14] , \Mem[8][13] ,
         \Mem[8][12] , \Mem[8][11] , \Mem[8][10] , \Mem[8][9] , \Mem[8][8] ,
         \Mem[8][7] , \Mem[8][6] , \Mem[8][5] , \Mem[8][4] , \Mem[8][3] ,
         \Mem[8][2] , \Mem[8][1] , \Mem[8][0] , \Mem[7][31] , \Mem[7][30] ,
         \Mem[7][29] , \Mem[7][28] , \Mem[7][27] , \Mem[7][26] , \Mem[7][25] ,
         \Mem[7][24] , \Mem[7][23] , \Mem[7][22] , \Mem[7][21] , \Mem[7][20] ,
         \Mem[7][19] , \Mem[7][18] , \Mem[7][17] , \Mem[7][16] , \Mem[7][15] ,
         \Mem[7][14] , \Mem[7][13] , \Mem[7][12] , \Mem[7][11] , \Mem[7][10] ,
         \Mem[7][9] , \Mem[7][8] , \Mem[7][7] , \Mem[7][6] , \Mem[7][5] ,
         \Mem[7][4] , \Mem[7][3] , \Mem[7][2] , \Mem[7][1] , \Mem[7][0] ,
         \Mem[6][31] , \Mem[6][30] , \Mem[6][29] , \Mem[6][28] , \Mem[6][27] ,
         \Mem[6][26] , \Mem[6][25] , \Mem[6][24] , \Mem[6][23] , \Mem[6][22] ,
         \Mem[6][21] , \Mem[6][20] , \Mem[6][19] , \Mem[6][18] , \Mem[6][17] ,
         \Mem[6][16] , \Mem[6][15] , \Mem[6][14] , \Mem[6][13] , \Mem[6][12] ,
         \Mem[6][11] , \Mem[6][10] , \Mem[6][9] , \Mem[6][8] , \Mem[6][7] ,
         \Mem[6][6] , \Mem[6][5] , \Mem[6][4] , \Mem[6][3] , \Mem[6][2] ,
         \Mem[6][1] , \Mem[6][0] , \Mem[5][31] , \Mem[5][30] , \Mem[5][29] ,
         \Mem[5][28] , \Mem[5][27] , \Mem[5][26] , \Mem[5][25] , \Mem[5][24] ,
         \Mem[5][23] , \Mem[5][22] , \Mem[5][21] , \Mem[5][20] , \Mem[5][19] ,
         \Mem[5][18] , \Mem[5][17] , \Mem[5][16] , \Mem[5][15] , \Mem[5][14] ,
         \Mem[5][13] , \Mem[5][12] , \Mem[5][11] , \Mem[5][10] , \Mem[5][9] ,
         \Mem[5][8] , \Mem[5][7] , \Mem[5][6] , \Mem[5][5] , \Mem[5][4] ,
         \Mem[5][3] , \Mem[5][2] , \Mem[5][1] , \Mem[5][0] , \Mem[4][31] ,
         \Mem[4][30] , \Mem[4][29] , \Mem[4][28] , \Mem[4][27] , \Mem[4][26] ,
         \Mem[4][25] , \Mem[4][24] , \Mem[4][23] , \Mem[4][22] , \Mem[4][21] ,
         \Mem[4][20] , \Mem[4][19] , \Mem[4][18] , \Mem[4][17] , \Mem[4][16] ,
         \Mem[4][15] , \Mem[4][14] , \Mem[4][13] , \Mem[4][12] , \Mem[4][11] ,
         \Mem[4][10] , \Mem[4][9] , \Mem[4][8] , \Mem[4][7] , \Mem[4][6] ,
         \Mem[4][5] , \Mem[4][4] , \Mem[4][3] , \Mem[4][2] , \Mem[4][1] ,
         \Mem[4][0] , \Mem[3][31] , \Mem[3][30] , \Mem[3][29] , \Mem[3][28] ,
         \Mem[3][27] , \Mem[3][26] , \Mem[3][25] , \Mem[3][24] , \Mem[3][23] ,
         \Mem[3][22] , \Mem[3][21] , \Mem[3][20] , \Mem[3][19] , \Mem[3][18] ,
         \Mem[3][17] , \Mem[3][16] , \Mem[3][15] , \Mem[3][14] , \Mem[3][13] ,
         \Mem[3][12] , \Mem[3][11] , \Mem[3][10] , \Mem[3][9] , \Mem[3][8] ,
         \Mem[3][7] , \Mem[3][6] , \Mem[3][5] , \Mem[3][4] , \Mem[3][3] ,
         \Mem[3][2] , \Mem[3][1] , \Mem[3][0] , \Mem[2][31] , \Mem[2][30] ,
         \Mem[2][29] , \Mem[2][28] , \Mem[2][27] , \Mem[2][26] , \Mem[2][25] ,
         \Mem[2][24] , \Mem[2][23] , \Mem[2][22] , \Mem[2][21] , \Mem[2][20] ,
         \Mem[2][19] , \Mem[2][18] , \Mem[2][17] , \Mem[2][16] , \Mem[2][15] ,
         \Mem[2][14] , \Mem[2][13] , \Mem[2][12] , \Mem[2][11] , \Mem[2][10] ,
         \Mem[2][9] , \Mem[2][8] , \Mem[2][7] , \Mem[2][6] , \Mem[2][5] ,
         \Mem[2][4] , \Mem[2][3] , \Mem[2][2] , \Mem[2][1] , \Mem[2][0] ,
         \Mem[1][31] , \Mem[1][30] , \Mem[1][29] , \Mem[1][28] , \Mem[1][27] ,
         \Mem[1][26] , \Mem[1][25] , \Mem[1][24] , \Mem[1][23] , \Mem[1][22] ,
         \Mem[1][21] , \Mem[1][20] , \Mem[1][19] , \Mem[1][18] , \Mem[1][17] ,
         \Mem[1][16] , \Mem[1][15] , \Mem[1][14] , \Mem[1][13] , \Mem[1][12] ,
         \Mem[1][11] , \Mem[1][10] , \Mem[1][9] , \Mem[1][8] , \Mem[1][7] ,
         \Mem[1][6] , \Mem[1][5] , \Mem[1][4] , \Mem[1][3] , \Mem[1][2] ,
         \Mem[1][1] , \Mem[1][0] , \Mem[0][31] , \Mem[0][30] , \Mem[0][29] ,
         \Mem[0][28] , \Mem[0][27] , \Mem[0][26] , \Mem[0][25] , \Mem[0][24] ,
         \Mem[0][23] , \Mem[0][22] , \Mem[0][21] , \Mem[0][20] , \Mem[0][19] ,
         \Mem[0][18] , \Mem[0][17] , \Mem[0][16] , \Mem[0][15] , \Mem[0][14] ,
         \Mem[0][13] , \Mem[0][12] , \Mem[0][11] , \Mem[0][10] , \Mem[0][9] ,
         \Mem[0][8] , \Mem[0][7] , \Mem[0][6] , \Mem[0][5] , \Mem[0][4] ,
         \Mem[0][3] , \Mem[0][2] , \Mem[0][1] , \Mem[0][0] , N81, N82, N83,
         N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97,
         N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109,
         N110, N111, N112, n1, n3, n5, n7, n9, n11, n13, n15, n17, n19, n21,
         n23, n25, n27, n28, n30, n32, n34, n36, n38, n40, n42, n44, n46, n48,
         n50, n52, n54, n56, n58, n60, n62, n64, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1957, n1958,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2219, n2220, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n80, n81, n115, n116, n150, n184,
         n218, n252, n286, n320, n356, n390, n623, n657, n923, n1190, n1456,
         n1722, n1956, n1959, n2025, n2026, n2027, n2218, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027;
  assign N10 = ADDR_RD[0];
  assign N11 = ADDR_RD[1];
  assign N12 = ADDR_RD[2];
  assign N13 = ADDR_RD[3];
  assign N14 = ADDR_RD[4];
  assign N15 = ADDR_RD[5];

  DFFPOSX1 \Mem_reg[63][31]  ( .D(n4333), .CLK(clk), .Q(\Mem[63][31] ) );
  DFFPOSX1 \Mem_reg[63][30]  ( .D(n4332), .CLK(clk), .Q(\Mem[63][30] ) );
  DFFPOSX1 \Mem_reg[63][29]  ( .D(n4331), .CLK(clk), .Q(\Mem[63][29] ) );
  DFFPOSX1 \Mem_reg[63][28]  ( .D(n4330), .CLK(clk), .Q(\Mem[63][28] ) );
  DFFPOSX1 \Mem_reg[63][27]  ( .D(n4329), .CLK(clk), .Q(\Mem[63][27] ) );
  DFFPOSX1 \Mem_reg[63][26]  ( .D(n4328), .CLK(clk), .Q(\Mem[63][26] ) );
  DFFPOSX1 \Mem_reg[63][25]  ( .D(n4327), .CLK(clk), .Q(\Mem[63][25] ) );
  DFFPOSX1 \Mem_reg[63][24]  ( .D(n4326), .CLK(clk), .Q(\Mem[63][24] ) );
  DFFPOSX1 \Mem_reg[63][23]  ( .D(n4325), .CLK(clk), .Q(\Mem[63][23] ) );
  DFFPOSX1 \Mem_reg[63][22]  ( .D(n4324), .CLK(clk), .Q(\Mem[63][22] ) );
  DFFPOSX1 \Mem_reg[63][21]  ( .D(n4323), .CLK(clk), .Q(\Mem[63][21] ) );
  DFFPOSX1 \Mem_reg[63][20]  ( .D(n4322), .CLK(clk), .Q(\Mem[63][20] ) );
  DFFPOSX1 \Mem_reg[63][19]  ( .D(n4321), .CLK(clk), .Q(\Mem[63][19] ) );
  DFFPOSX1 \Mem_reg[63][18]  ( .D(n4320), .CLK(clk), .Q(\Mem[63][18] ) );
  DFFPOSX1 \Mem_reg[63][17]  ( .D(n4319), .CLK(clk), .Q(\Mem[63][17] ) );
  DFFPOSX1 \Mem_reg[63][16]  ( .D(n4318), .CLK(clk), .Q(\Mem[63][16] ) );
  DFFPOSX1 \Mem_reg[63][15]  ( .D(n4317), .CLK(clk), .Q(\Mem[63][15] ) );
  DFFPOSX1 \Mem_reg[63][14]  ( .D(n4316), .CLK(clk), .Q(\Mem[63][14] ) );
  DFFPOSX1 \Mem_reg[63][13]  ( .D(n4315), .CLK(clk), .Q(\Mem[63][13] ) );
  DFFPOSX1 \Mem_reg[63][12]  ( .D(n4314), .CLK(clk), .Q(\Mem[63][12] ) );
  DFFPOSX1 \Mem_reg[63][11]  ( .D(n4313), .CLK(clk), .Q(\Mem[63][11] ) );
  DFFPOSX1 \Mem_reg[63][10]  ( .D(n4312), .CLK(clk), .Q(\Mem[63][10] ) );
  DFFPOSX1 \Mem_reg[63][9]  ( .D(n4311), .CLK(clk), .Q(\Mem[63][9] ) );
  DFFPOSX1 \Mem_reg[63][8]  ( .D(n4310), .CLK(clk), .Q(\Mem[63][8] ) );
  DFFPOSX1 \Mem_reg[63][7]  ( .D(n4309), .CLK(clk), .Q(\Mem[63][7] ) );
  DFFPOSX1 \Mem_reg[63][6]  ( .D(n4308), .CLK(clk), .Q(\Mem[63][6] ) );
  DFFPOSX1 \Mem_reg[63][5]  ( .D(n4307), .CLK(clk), .Q(\Mem[63][5] ) );
  DFFPOSX1 \Mem_reg[63][4]  ( .D(n4306), .CLK(clk), .Q(\Mem[63][4] ) );
  DFFPOSX1 \Mem_reg[63][3]  ( .D(n4305), .CLK(clk), .Q(\Mem[63][3] ) );
  DFFPOSX1 \Mem_reg[63][2]  ( .D(n4304), .CLK(clk), .Q(\Mem[63][2] ) );
  DFFPOSX1 \Mem_reg[63][1]  ( .D(n4303), .CLK(clk), .Q(\Mem[63][1] ) );
  DFFPOSX1 \Mem_reg[63][0]  ( .D(n4302), .CLK(clk), .Q(\Mem[63][0] ) );
  DFFPOSX1 \Mem_reg[62][31]  ( .D(n4301), .CLK(clk), .Q(\Mem[62][31] ) );
  DFFPOSX1 \Mem_reg[62][30]  ( .D(n4300), .CLK(clk), .Q(\Mem[62][30] ) );
  DFFPOSX1 \Mem_reg[62][29]  ( .D(n4299), .CLK(clk), .Q(\Mem[62][29] ) );
  DFFPOSX1 \Mem_reg[62][28]  ( .D(n4298), .CLK(clk), .Q(\Mem[62][28] ) );
  DFFPOSX1 \Mem_reg[62][27]  ( .D(n4297), .CLK(clk), .Q(\Mem[62][27] ) );
  DFFPOSX1 \Mem_reg[62][26]  ( .D(n4296), .CLK(clk), .Q(\Mem[62][26] ) );
  DFFPOSX1 \Mem_reg[62][25]  ( .D(n4295), .CLK(clk), .Q(\Mem[62][25] ) );
  DFFPOSX1 \Mem_reg[62][24]  ( .D(n4294), .CLK(clk), .Q(\Mem[62][24] ) );
  DFFPOSX1 \Mem_reg[62][23]  ( .D(n4293), .CLK(clk), .Q(\Mem[62][23] ) );
  DFFPOSX1 \Mem_reg[62][22]  ( .D(n4292), .CLK(clk), .Q(\Mem[62][22] ) );
  DFFPOSX1 \Mem_reg[62][21]  ( .D(n4291), .CLK(clk), .Q(\Mem[62][21] ) );
  DFFPOSX1 \Mem_reg[62][20]  ( .D(n4290), .CLK(clk), .Q(\Mem[62][20] ) );
  DFFPOSX1 \Mem_reg[62][19]  ( .D(n4289), .CLK(clk), .Q(\Mem[62][19] ) );
  DFFPOSX1 \Mem_reg[62][18]  ( .D(n4288), .CLK(clk), .Q(\Mem[62][18] ) );
  DFFPOSX1 \Mem_reg[62][17]  ( .D(n4287), .CLK(clk), .Q(\Mem[62][17] ) );
  DFFPOSX1 \Mem_reg[62][16]  ( .D(n4286), .CLK(clk), .Q(\Mem[62][16] ) );
  DFFPOSX1 \Mem_reg[62][15]  ( .D(n4285), .CLK(clk), .Q(\Mem[62][15] ) );
  DFFPOSX1 \Mem_reg[62][14]  ( .D(n4284), .CLK(clk), .Q(\Mem[62][14] ) );
  DFFPOSX1 \Mem_reg[62][13]  ( .D(n4283), .CLK(clk), .Q(\Mem[62][13] ) );
  DFFPOSX1 \Mem_reg[62][12]  ( .D(n4282), .CLK(clk), .Q(\Mem[62][12] ) );
  DFFPOSX1 \Mem_reg[62][11]  ( .D(n4281), .CLK(clk), .Q(\Mem[62][11] ) );
  DFFPOSX1 \Mem_reg[62][10]  ( .D(n4280), .CLK(clk), .Q(\Mem[62][10] ) );
  DFFPOSX1 \Mem_reg[62][9]  ( .D(n4279), .CLK(clk), .Q(\Mem[62][9] ) );
  DFFPOSX1 \Mem_reg[62][8]  ( .D(n4278), .CLK(clk), .Q(\Mem[62][8] ) );
  DFFPOSX1 \Mem_reg[62][7]  ( .D(n4277), .CLK(clk), .Q(\Mem[62][7] ) );
  DFFPOSX1 \Mem_reg[62][6]  ( .D(n4276), .CLK(clk), .Q(\Mem[62][6] ) );
  DFFPOSX1 \Mem_reg[62][5]  ( .D(n4275), .CLK(clk), .Q(\Mem[62][5] ) );
  DFFPOSX1 \Mem_reg[62][4]  ( .D(n4274), .CLK(clk), .Q(\Mem[62][4] ) );
  DFFPOSX1 \Mem_reg[62][3]  ( .D(n4273), .CLK(clk), .Q(\Mem[62][3] ) );
  DFFPOSX1 \Mem_reg[62][2]  ( .D(n4272), .CLK(clk), .Q(\Mem[62][2] ) );
  DFFPOSX1 \Mem_reg[62][1]  ( .D(n4271), .CLK(clk), .Q(\Mem[62][1] ) );
  DFFPOSX1 \Mem_reg[62][0]  ( .D(n4270), .CLK(clk), .Q(\Mem[62][0] ) );
  DFFPOSX1 \Mem_reg[61][31]  ( .D(n4269), .CLK(clk), .Q(\Mem[61][31] ) );
  DFFPOSX1 \Mem_reg[61][30]  ( .D(n4268), .CLK(clk), .Q(\Mem[61][30] ) );
  DFFPOSX1 \Mem_reg[61][29]  ( .D(n4267), .CLK(clk), .Q(\Mem[61][29] ) );
  DFFPOSX1 \Mem_reg[61][28]  ( .D(n4266), .CLK(clk), .Q(\Mem[61][28] ) );
  DFFPOSX1 \Mem_reg[61][27]  ( .D(n4265), .CLK(clk), .Q(\Mem[61][27] ) );
  DFFPOSX1 \Mem_reg[61][26]  ( .D(n4264), .CLK(clk), .Q(\Mem[61][26] ) );
  DFFPOSX1 \Mem_reg[61][25]  ( .D(n4263), .CLK(clk), .Q(\Mem[61][25] ) );
  DFFPOSX1 \Mem_reg[61][24]  ( .D(n4262), .CLK(clk), .Q(\Mem[61][24] ) );
  DFFPOSX1 \Mem_reg[61][23]  ( .D(n4261), .CLK(clk), .Q(\Mem[61][23] ) );
  DFFPOSX1 \Mem_reg[61][22]  ( .D(n4260), .CLK(clk), .Q(\Mem[61][22] ) );
  DFFPOSX1 \Mem_reg[61][21]  ( .D(n4259), .CLK(clk), .Q(\Mem[61][21] ) );
  DFFPOSX1 \Mem_reg[61][20]  ( .D(n4258), .CLK(clk), .Q(\Mem[61][20] ) );
  DFFPOSX1 \Mem_reg[61][19]  ( .D(n4257), .CLK(clk), .Q(\Mem[61][19] ) );
  DFFPOSX1 \Mem_reg[61][18]  ( .D(n4256), .CLK(clk), .Q(\Mem[61][18] ) );
  DFFPOSX1 \Mem_reg[61][17]  ( .D(n4255), .CLK(clk), .Q(\Mem[61][17] ) );
  DFFPOSX1 \Mem_reg[61][16]  ( .D(n4254), .CLK(clk), .Q(\Mem[61][16] ) );
  DFFPOSX1 \Mem_reg[61][15]  ( .D(n4253), .CLK(clk), .Q(\Mem[61][15] ) );
  DFFPOSX1 \Mem_reg[61][14]  ( .D(n4252), .CLK(clk), .Q(\Mem[61][14] ) );
  DFFPOSX1 \Mem_reg[61][13]  ( .D(n4251), .CLK(clk), .Q(\Mem[61][13] ) );
  DFFPOSX1 \Mem_reg[61][12]  ( .D(n4250), .CLK(clk), .Q(\Mem[61][12] ) );
  DFFPOSX1 \Mem_reg[61][11]  ( .D(n4249), .CLK(clk), .Q(\Mem[61][11] ) );
  DFFPOSX1 \Mem_reg[61][10]  ( .D(n4248), .CLK(clk), .Q(\Mem[61][10] ) );
  DFFPOSX1 \Mem_reg[61][9]  ( .D(n4247), .CLK(clk), .Q(\Mem[61][9] ) );
  DFFPOSX1 \Mem_reg[61][8]  ( .D(n4246), .CLK(clk), .Q(\Mem[61][8] ) );
  DFFPOSX1 \Mem_reg[61][7]  ( .D(n4245), .CLK(clk), .Q(\Mem[61][7] ) );
  DFFPOSX1 \Mem_reg[61][6]  ( .D(n4244), .CLK(clk), .Q(\Mem[61][6] ) );
  DFFPOSX1 \Mem_reg[61][5]  ( .D(n4243), .CLK(clk), .Q(\Mem[61][5] ) );
  DFFPOSX1 \Mem_reg[61][4]  ( .D(n4242), .CLK(clk), .Q(\Mem[61][4] ) );
  DFFPOSX1 \Mem_reg[61][3]  ( .D(n4241), .CLK(clk), .Q(\Mem[61][3] ) );
  DFFPOSX1 \Mem_reg[61][2]  ( .D(n4240), .CLK(clk), .Q(\Mem[61][2] ) );
  DFFPOSX1 \Mem_reg[61][1]  ( .D(n4239), .CLK(clk), .Q(\Mem[61][1] ) );
  DFFPOSX1 \Mem_reg[61][0]  ( .D(n4238), .CLK(clk), .Q(\Mem[61][0] ) );
  DFFPOSX1 \Mem_reg[60][31]  ( .D(n4237), .CLK(clk), .Q(\Mem[60][31] ) );
  DFFPOSX1 \Mem_reg[60][30]  ( .D(n4236), .CLK(clk), .Q(\Mem[60][30] ) );
  DFFPOSX1 \Mem_reg[60][29]  ( .D(n4235), .CLK(clk), .Q(\Mem[60][29] ) );
  DFFPOSX1 \Mem_reg[60][28]  ( .D(n4234), .CLK(clk), .Q(\Mem[60][28] ) );
  DFFPOSX1 \Mem_reg[60][27]  ( .D(n4233), .CLK(clk), .Q(\Mem[60][27] ) );
  DFFPOSX1 \Mem_reg[60][26]  ( .D(n4232), .CLK(clk), .Q(\Mem[60][26] ) );
  DFFPOSX1 \Mem_reg[60][25]  ( .D(n4231), .CLK(clk), .Q(\Mem[60][25] ) );
  DFFPOSX1 \Mem_reg[60][24]  ( .D(n4230), .CLK(clk), .Q(\Mem[60][24] ) );
  DFFPOSX1 \Mem_reg[60][23]  ( .D(n4229), .CLK(clk), .Q(\Mem[60][23] ) );
  DFFPOSX1 \Mem_reg[60][22]  ( .D(n4228), .CLK(clk), .Q(\Mem[60][22] ) );
  DFFPOSX1 \Mem_reg[60][21]  ( .D(n4227), .CLK(clk), .Q(\Mem[60][21] ) );
  DFFPOSX1 \Mem_reg[60][20]  ( .D(n4226), .CLK(clk), .Q(\Mem[60][20] ) );
  DFFPOSX1 \Mem_reg[60][19]  ( .D(n4225), .CLK(clk), .Q(\Mem[60][19] ) );
  DFFPOSX1 \Mem_reg[60][18]  ( .D(n4224), .CLK(clk), .Q(\Mem[60][18] ) );
  DFFPOSX1 \Mem_reg[60][17]  ( .D(n4223), .CLK(clk), .Q(\Mem[60][17] ) );
  DFFPOSX1 \Mem_reg[60][16]  ( .D(n4222), .CLK(clk), .Q(\Mem[60][16] ) );
  DFFPOSX1 \Mem_reg[60][15]  ( .D(n4221), .CLK(clk), .Q(\Mem[60][15] ) );
  DFFPOSX1 \Mem_reg[60][14]  ( .D(n4220), .CLK(clk), .Q(\Mem[60][14] ) );
  DFFPOSX1 \Mem_reg[60][13]  ( .D(n4219), .CLK(clk), .Q(\Mem[60][13] ) );
  DFFPOSX1 \Mem_reg[60][12]  ( .D(n4218), .CLK(clk), .Q(\Mem[60][12] ) );
  DFFPOSX1 \Mem_reg[60][11]  ( .D(n4217), .CLK(clk), .Q(\Mem[60][11] ) );
  DFFPOSX1 \Mem_reg[60][10]  ( .D(n4216), .CLK(clk), .Q(\Mem[60][10] ) );
  DFFPOSX1 \Mem_reg[60][9]  ( .D(n4215), .CLK(clk), .Q(\Mem[60][9] ) );
  DFFPOSX1 \Mem_reg[60][8]  ( .D(n4214), .CLK(clk), .Q(\Mem[60][8] ) );
  DFFPOSX1 \Mem_reg[60][7]  ( .D(n4213), .CLK(clk), .Q(\Mem[60][7] ) );
  DFFPOSX1 \Mem_reg[60][6]  ( .D(n4212), .CLK(clk), .Q(\Mem[60][6] ) );
  DFFPOSX1 \Mem_reg[60][5]  ( .D(n4211), .CLK(clk), .Q(\Mem[60][5] ) );
  DFFPOSX1 \Mem_reg[60][4]  ( .D(n4210), .CLK(clk), .Q(\Mem[60][4] ) );
  DFFPOSX1 \Mem_reg[60][3]  ( .D(n4209), .CLK(clk), .Q(\Mem[60][3] ) );
  DFFPOSX1 \Mem_reg[60][2]  ( .D(n4208), .CLK(clk), .Q(\Mem[60][2] ) );
  DFFPOSX1 \Mem_reg[60][1]  ( .D(n4207), .CLK(clk), .Q(\Mem[60][1] ) );
  DFFPOSX1 \Mem_reg[60][0]  ( .D(n4206), .CLK(clk), .Q(\Mem[60][0] ) );
  DFFPOSX1 \Mem_reg[59][31]  ( .D(n4205), .CLK(clk), .Q(\Mem[59][31] ) );
  DFFPOSX1 \Mem_reg[59][30]  ( .D(n4204), .CLK(clk), .Q(\Mem[59][30] ) );
  DFFPOSX1 \Mem_reg[59][29]  ( .D(n4203), .CLK(clk), .Q(\Mem[59][29] ) );
  DFFPOSX1 \Mem_reg[59][28]  ( .D(n4202), .CLK(clk), .Q(\Mem[59][28] ) );
  DFFPOSX1 \Mem_reg[59][27]  ( .D(n4201), .CLK(clk), .Q(\Mem[59][27] ) );
  DFFPOSX1 \Mem_reg[59][26]  ( .D(n4200), .CLK(clk), .Q(\Mem[59][26] ) );
  DFFPOSX1 \Mem_reg[59][25]  ( .D(n4199), .CLK(clk), .Q(\Mem[59][25] ) );
  DFFPOSX1 \Mem_reg[59][24]  ( .D(n4198), .CLK(clk), .Q(\Mem[59][24] ) );
  DFFPOSX1 \Mem_reg[59][23]  ( .D(n4197), .CLK(clk), .Q(\Mem[59][23] ) );
  DFFPOSX1 \Mem_reg[59][22]  ( .D(n4196), .CLK(clk), .Q(\Mem[59][22] ) );
  DFFPOSX1 \Mem_reg[59][21]  ( .D(n4195), .CLK(clk), .Q(\Mem[59][21] ) );
  DFFPOSX1 \Mem_reg[59][20]  ( .D(n4194), .CLK(clk), .Q(\Mem[59][20] ) );
  DFFPOSX1 \Mem_reg[59][19]  ( .D(n4193), .CLK(clk), .Q(\Mem[59][19] ) );
  DFFPOSX1 \Mem_reg[59][18]  ( .D(n4192), .CLK(clk), .Q(\Mem[59][18] ) );
  DFFPOSX1 \Mem_reg[59][17]  ( .D(n4191), .CLK(clk), .Q(\Mem[59][17] ) );
  DFFPOSX1 \Mem_reg[59][16]  ( .D(n4190), .CLK(clk), .Q(\Mem[59][16] ) );
  DFFPOSX1 \Mem_reg[59][15]  ( .D(n4189), .CLK(clk), .Q(\Mem[59][15] ) );
  DFFPOSX1 \Mem_reg[59][14]  ( .D(n4188), .CLK(clk), .Q(\Mem[59][14] ) );
  DFFPOSX1 \Mem_reg[59][13]  ( .D(n4187), .CLK(clk), .Q(\Mem[59][13] ) );
  DFFPOSX1 \Mem_reg[59][12]  ( .D(n4186), .CLK(clk), .Q(\Mem[59][12] ) );
  DFFPOSX1 \Mem_reg[59][11]  ( .D(n4185), .CLK(clk), .Q(\Mem[59][11] ) );
  DFFPOSX1 \Mem_reg[59][10]  ( .D(n4184), .CLK(clk), .Q(\Mem[59][10] ) );
  DFFPOSX1 \Mem_reg[59][9]  ( .D(n4183), .CLK(clk), .Q(\Mem[59][9] ) );
  DFFPOSX1 \Mem_reg[59][8]  ( .D(n4182), .CLK(clk), .Q(\Mem[59][8] ) );
  DFFPOSX1 \Mem_reg[59][7]  ( .D(n4181), .CLK(clk), .Q(\Mem[59][7] ) );
  DFFPOSX1 \Mem_reg[59][6]  ( .D(n4180), .CLK(clk), .Q(\Mem[59][6] ) );
  DFFPOSX1 \Mem_reg[59][5]  ( .D(n4179), .CLK(clk), .Q(\Mem[59][5] ) );
  DFFPOSX1 \Mem_reg[59][4]  ( .D(n4178), .CLK(clk), .Q(\Mem[59][4] ) );
  DFFPOSX1 \Mem_reg[59][3]  ( .D(n4177), .CLK(clk), .Q(\Mem[59][3] ) );
  DFFPOSX1 \Mem_reg[59][2]  ( .D(n4176), .CLK(clk), .Q(\Mem[59][2] ) );
  DFFPOSX1 \Mem_reg[59][1]  ( .D(n4175), .CLK(clk), .Q(\Mem[59][1] ) );
  DFFPOSX1 \Mem_reg[59][0]  ( .D(n4174), .CLK(clk), .Q(\Mem[59][0] ) );
  DFFPOSX1 \Mem_reg[58][31]  ( .D(n4173), .CLK(clk), .Q(\Mem[58][31] ) );
  DFFPOSX1 \Mem_reg[58][30]  ( .D(n4172), .CLK(clk), .Q(\Mem[58][30] ) );
  DFFPOSX1 \Mem_reg[58][29]  ( .D(n4171), .CLK(clk), .Q(\Mem[58][29] ) );
  DFFPOSX1 \Mem_reg[58][28]  ( .D(n4170), .CLK(clk), .Q(\Mem[58][28] ) );
  DFFPOSX1 \Mem_reg[58][27]  ( .D(n4169), .CLK(clk), .Q(\Mem[58][27] ) );
  DFFPOSX1 \Mem_reg[58][26]  ( .D(n4168), .CLK(clk), .Q(\Mem[58][26] ) );
  DFFPOSX1 \Mem_reg[58][25]  ( .D(n4167), .CLK(clk), .Q(\Mem[58][25] ) );
  DFFPOSX1 \Mem_reg[58][24]  ( .D(n4166), .CLK(clk), .Q(\Mem[58][24] ) );
  DFFPOSX1 \Mem_reg[58][23]  ( .D(n4165), .CLK(clk), .Q(\Mem[58][23] ) );
  DFFPOSX1 \Mem_reg[58][22]  ( .D(n4164), .CLK(clk), .Q(\Mem[58][22] ) );
  DFFPOSX1 \Mem_reg[58][21]  ( .D(n4163), .CLK(clk), .Q(\Mem[58][21] ) );
  DFFPOSX1 \Mem_reg[58][20]  ( .D(n4162), .CLK(clk), .Q(\Mem[58][20] ) );
  DFFPOSX1 \Mem_reg[58][19]  ( .D(n4161), .CLK(clk), .Q(\Mem[58][19] ) );
  DFFPOSX1 \Mem_reg[58][18]  ( .D(n4160), .CLK(clk), .Q(\Mem[58][18] ) );
  DFFPOSX1 \Mem_reg[58][17]  ( .D(n4159), .CLK(clk), .Q(\Mem[58][17] ) );
  DFFPOSX1 \Mem_reg[58][16]  ( .D(n4158), .CLK(clk), .Q(\Mem[58][16] ) );
  DFFPOSX1 \Mem_reg[58][15]  ( .D(n4157), .CLK(clk), .Q(\Mem[58][15] ) );
  DFFPOSX1 \Mem_reg[58][14]  ( .D(n4156), .CLK(clk), .Q(\Mem[58][14] ) );
  DFFPOSX1 \Mem_reg[58][13]  ( .D(n4155), .CLK(clk), .Q(\Mem[58][13] ) );
  DFFPOSX1 \Mem_reg[58][12]  ( .D(n4154), .CLK(clk), .Q(\Mem[58][12] ) );
  DFFPOSX1 \Mem_reg[58][11]  ( .D(n4153), .CLK(clk), .Q(\Mem[58][11] ) );
  DFFPOSX1 \Mem_reg[58][10]  ( .D(n4152), .CLK(clk), .Q(\Mem[58][10] ) );
  DFFPOSX1 \Mem_reg[58][9]  ( .D(n4151), .CLK(clk), .Q(\Mem[58][9] ) );
  DFFPOSX1 \Mem_reg[58][8]  ( .D(n4150), .CLK(clk), .Q(\Mem[58][8] ) );
  DFFPOSX1 \Mem_reg[58][7]  ( .D(n4149), .CLK(clk), .Q(\Mem[58][7] ) );
  DFFPOSX1 \Mem_reg[58][6]  ( .D(n4148), .CLK(clk), .Q(\Mem[58][6] ) );
  DFFPOSX1 \Mem_reg[58][5]  ( .D(n4147), .CLK(clk), .Q(\Mem[58][5] ) );
  DFFPOSX1 \Mem_reg[58][4]  ( .D(n4146), .CLK(clk), .Q(\Mem[58][4] ) );
  DFFPOSX1 \Mem_reg[58][3]  ( .D(n4145), .CLK(clk), .Q(\Mem[58][3] ) );
  DFFPOSX1 \Mem_reg[58][2]  ( .D(n4144), .CLK(clk), .Q(\Mem[58][2] ) );
  DFFPOSX1 \Mem_reg[58][1]  ( .D(n4143), .CLK(clk), .Q(\Mem[58][1] ) );
  DFFPOSX1 \Mem_reg[58][0]  ( .D(n4142), .CLK(clk), .Q(\Mem[58][0] ) );
  DFFPOSX1 \Mem_reg[57][31]  ( .D(n4141), .CLK(clk), .Q(\Mem[57][31] ) );
  DFFPOSX1 \Mem_reg[57][30]  ( .D(n4140), .CLK(clk), .Q(\Mem[57][30] ) );
  DFFPOSX1 \Mem_reg[57][29]  ( .D(n4139), .CLK(clk), .Q(\Mem[57][29] ) );
  DFFPOSX1 \Mem_reg[57][28]  ( .D(n4138), .CLK(clk), .Q(\Mem[57][28] ) );
  DFFPOSX1 \Mem_reg[57][27]  ( .D(n4137), .CLK(clk), .Q(\Mem[57][27] ) );
  DFFPOSX1 \Mem_reg[57][26]  ( .D(n4136), .CLK(clk), .Q(\Mem[57][26] ) );
  DFFPOSX1 \Mem_reg[57][25]  ( .D(n4135), .CLK(clk), .Q(\Mem[57][25] ) );
  DFFPOSX1 \Mem_reg[57][24]  ( .D(n4134), .CLK(clk), .Q(\Mem[57][24] ) );
  DFFPOSX1 \Mem_reg[57][23]  ( .D(n4133), .CLK(clk), .Q(\Mem[57][23] ) );
  DFFPOSX1 \Mem_reg[57][22]  ( .D(n4132), .CLK(clk), .Q(\Mem[57][22] ) );
  DFFPOSX1 \Mem_reg[57][21]  ( .D(n4131), .CLK(clk), .Q(\Mem[57][21] ) );
  DFFPOSX1 \Mem_reg[57][20]  ( .D(n4130), .CLK(clk), .Q(\Mem[57][20] ) );
  DFFPOSX1 \Mem_reg[57][19]  ( .D(n4129), .CLK(clk), .Q(\Mem[57][19] ) );
  DFFPOSX1 \Mem_reg[57][18]  ( .D(n4128), .CLK(clk), .Q(\Mem[57][18] ) );
  DFFPOSX1 \Mem_reg[57][17]  ( .D(n4127), .CLK(clk), .Q(\Mem[57][17] ) );
  DFFPOSX1 \Mem_reg[57][16]  ( .D(n4126), .CLK(clk), .Q(\Mem[57][16] ) );
  DFFPOSX1 \Mem_reg[57][15]  ( .D(n4125), .CLK(clk), .Q(\Mem[57][15] ) );
  DFFPOSX1 \Mem_reg[57][14]  ( .D(n4124), .CLK(clk), .Q(\Mem[57][14] ) );
  DFFPOSX1 \Mem_reg[57][13]  ( .D(n4123), .CLK(clk), .Q(\Mem[57][13] ) );
  DFFPOSX1 \Mem_reg[57][12]  ( .D(n4122), .CLK(clk), .Q(\Mem[57][12] ) );
  DFFPOSX1 \Mem_reg[57][11]  ( .D(n4121), .CLK(clk), .Q(\Mem[57][11] ) );
  DFFPOSX1 \Mem_reg[57][10]  ( .D(n4120), .CLK(clk), .Q(\Mem[57][10] ) );
  DFFPOSX1 \Mem_reg[57][9]  ( .D(n4119), .CLK(clk), .Q(\Mem[57][9] ) );
  DFFPOSX1 \Mem_reg[57][8]  ( .D(n4118), .CLK(clk), .Q(\Mem[57][8] ) );
  DFFPOSX1 \Mem_reg[57][7]  ( .D(n4117), .CLK(clk), .Q(\Mem[57][7] ) );
  DFFPOSX1 \Mem_reg[57][6]  ( .D(n4116), .CLK(clk), .Q(\Mem[57][6] ) );
  DFFPOSX1 \Mem_reg[57][5]  ( .D(n4115), .CLK(clk), .Q(\Mem[57][5] ) );
  DFFPOSX1 \Mem_reg[57][4]  ( .D(n4114), .CLK(clk), .Q(\Mem[57][4] ) );
  DFFPOSX1 \Mem_reg[57][3]  ( .D(n4113), .CLK(clk), .Q(\Mem[57][3] ) );
  DFFPOSX1 \Mem_reg[57][2]  ( .D(n4112), .CLK(clk), .Q(\Mem[57][2] ) );
  DFFPOSX1 \Mem_reg[57][1]  ( .D(n4111), .CLK(clk), .Q(\Mem[57][1] ) );
  DFFPOSX1 \Mem_reg[57][0]  ( .D(n4110), .CLK(clk), .Q(\Mem[57][0] ) );
  DFFPOSX1 \Mem_reg[56][31]  ( .D(n4109), .CLK(clk), .Q(\Mem[56][31] ) );
  DFFPOSX1 \Mem_reg[56][30]  ( .D(n4108), .CLK(clk), .Q(\Mem[56][30] ) );
  DFFPOSX1 \Mem_reg[56][29]  ( .D(n4107), .CLK(clk), .Q(\Mem[56][29] ) );
  DFFPOSX1 \Mem_reg[56][28]  ( .D(n4106), .CLK(clk), .Q(\Mem[56][28] ) );
  DFFPOSX1 \Mem_reg[56][27]  ( .D(n4105), .CLK(clk), .Q(\Mem[56][27] ) );
  DFFPOSX1 \Mem_reg[56][26]  ( .D(n4104), .CLK(clk), .Q(\Mem[56][26] ) );
  DFFPOSX1 \Mem_reg[56][25]  ( .D(n4103), .CLK(clk), .Q(\Mem[56][25] ) );
  DFFPOSX1 \Mem_reg[56][24]  ( .D(n4102), .CLK(clk), .Q(\Mem[56][24] ) );
  DFFPOSX1 \Mem_reg[56][23]  ( .D(n4101), .CLK(clk), .Q(\Mem[56][23] ) );
  DFFPOSX1 \Mem_reg[56][22]  ( .D(n4100), .CLK(clk), .Q(\Mem[56][22] ) );
  DFFPOSX1 \Mem_reg[56][21]  ( .D(n4099), .CLK(clk), .Q(\Mem[56][21] ) );
  DFFPOSX1 \Mem_reg[56][20]  ( .D(n4098), .CLK(clk), .Q(\Mem[56][20] ) );
  DFFPOSX1 \Mem_reg[56][19]  ( .D(n4097), .CLK(clk), .Q(\Mem[56][19] ) );
  DFFPOSX1 \Mem_reg[56][18]  ( .D(n4096), .CLK(clk), .Q(\Mem[56][18] ) );
  DFFPOSX1 \Mem_reg[56][17]  ( .D(n4095), .CLK(clk), .Q(\Mem[56][17] ) );
  DFFPOSX1 \Mem_reg[56][16]  ( .D(n4094), .CLK(clk), .Q(\Mem[56][16] ) );
  DFFPOSX1 \Mem_reg[56][15]  ( .D(n4093), .CLK(clk), .Q(\Mem[56][15] ) );
  DFFPOSX1 \Mem_reg[56][14]  ( .D(n4092), .CLK(clk), .Q(\Mem[56][14] ) );
  DFFPOSX1 \Mem_reg[56][13]  ( .D(n4091), .CLK(clk), .Q(\Mem[56][13] ) );
  DFFPOSX1 \Mem_reg[56][12]  ( .D(n4090), .CLK(clk), .Q(\Mem[56][12] ) );
  DFFPOSX1 \Mem_reg[56][11]  ( .D(n4089), .CLK(clk), .Q(\Mem[56][11] ) );
  DFFPOSX1 \Mem_reg[56][10]  ( .D(n4088), .CLK(clk), .Q(\Mem[56][10] ) );
  DFFPOSX1 \Mem_reg[56][9]  ( .D(n4087), .CLK(clk), .Q(\Mem[56][9] ) );
  DFFPOSX1 \Mem_reg[56][8]  ( .D(n4086), .CLK(clk), .Q(\Mem[56][8] ) );
  DFFPOSX1 \Mem_reg[56][7]  ( .D(n4085), .CLK(clk), .Q(\Mem[56][7] ) );
  DFFPOSX1 \Mem_reg[56][6]  ( .D(n4084), .CLK(clk), .Q(\Mem[56][6] ) );
  DFFPOSX1 \Mem_reg[56][5]  ( .D(n4083), .CLK(clk), .Q(\Mem[56][5] ) );
  DFFPOSX1 \Mem_reg[56][4]  ( .D(n4082), .CLK(clk), .Q(\Mem[56][4] ) );
  DFFPOSX1 \Mem_reg[56][3]  ( .D(n4081), .CLK(clk), .Q(\Mem[56][3] ) );
  DFFPOSX1 \Mem_reg[56][2]  ( .D(n4080), .CLK(clk), .Q(\Mem[56][2] ) );
  DFFPOSX1 \Mem_reg[56][1]  ( .D(n4079), .CLK(clk), .Q(\Mem[56][1] ) );
  DFFPOSX1 \Mem_reg[56][0]  ( .D(n4078), .CLK(clk), .Q(\Mem[56][0] ) );
  DFFPOSX1 \Mem_reg[55][31]  ( .D(n4077), .CLK(clk), .Q(\Mem[55][31] ) );
  DFFPOSX1 \Mem_reg[55][30]  ( .D(n4076), .CLK(clk), .Q(\Mem[55][30] ) );
  DFFPOSX1 \Mem_reg[55][29]  ( .D(n4075), .CLK(clk), .Q(\Mem[55][29] ) );
  DFFPOSX1 \Mem_reg[55][28]  ( .D(n4074), .CLK(clk), .Q(\Mem[55][28] ) );
  DFFPOSX1 \Mem_reg[55][27]  ( .D(n4073), .CLK(clk), .Q(\Mem[55][27] ) );
  DFFPOSX1 \Mem_reg[55][26]  ( .D(n4072), .CLK(clk), .Q(\Mem[55][26] ) );
  DFFPOSX1 \Mem_reg[55][25]  ( .D(n4071), .CLK(clk), .Q(\Mem[55][25] ) );
  DFFPOSX1 \Mem_reg[55][24]  ( .D(n4070), .CLK(clk), .Q(\Mem[55][24] ) );
  DFFPOSX1 \Mem_reg[55][23]  ( .D(n4069), .CLK(clk), .Q(\Mem[55][23] ) );
  DFFPOSX1 \Mem_reg[55][22]  ( .D(n4068), .CLK(clk), .Q(\Mem[55][22] ) );
  DFFPOSX1 \Mem_reg[55][21]  ( .D(n4067), .CLK(clk), .Q(\Mem[55][21] ) );
  DFFPOSX1 \Mem_reg[55][20]  ( .D(n4066), .CLK(clk), .Q(\Mem[55][20] ) );
  DFFPOSX1 \Mem_reg[55][19]  ( .D(n4065), .CLK(clk), .Q(\Mem[55][19] ) );
  DFFPOSX1 \Mem_reg[55][18]  ( .D(n4064), .CLK(clk), .Q(\Mem[55][18] ) );
  DFFPOSX1 \Mem_reg[55][17]  ( .D(n4063), .CLK(clk), .Q(\Mem[55][17] ) );
  DFFPOSX1 \Mem_reg[55][16]  ( .D(n4062), .CLK(clk), .Q(\Mem[55][16] ) );
  DFFPOSX1 \Mem_reg[55][15]  ( .D(n4061), .CLK(clk), .Q(\Mem[55][15] ) );
  DFFPOSX1 \Mem_reg[55][14]  ( .D(n4060), .CLK(clk), .Q(\Mem[55][14] ) );
  DFFPOSX1 \Mem_reg[55][13]  ( .D(n4059), .CLK(clk), .Q(\Mem[55][13] ) );
  DFFPOSX1 \Mem_reg[55][12]  ( .D(n4058), .CLK(clk), .Q(\Mem[55][12] ) );
  DFFPOSX1 \Mem_reg[55][11]  ( .D(n4057), .CLK(clk), .Q(\Mem[55][11] ) );
  DFFPOSX1 \Mem_reg[55][10]  ( .D(n4056), .CLK(clk), .Q(\Mem[55][10] ) );
  DFFPOSX1 \Mem_reg[55][9]  ( .D(n4055), .CLK(clk), .Q(\Mem[55][9] ) );
  DFFPOSX1 \Mem_reg[55][8]  ( .D(n4054), .CLK(clk), .Q(\Mem[55][8] ) );
  DFFPOSX1 \Mem_reg[55][7]  ( .D(n4053), .CLK(clk), .Q(\Mem[55][7] ) );
  DFFPOSX1 \Mem_reg[55][6]  ( .D(n4052), .CLK(clk), .Q(\Mem[55][6] ) );
  DFFPOSX1 \Mem_reg[55][5]  ( .D(n4051), .CLK(clk), .Q(\Mem[55][5] ) );
  DFFPOSX1 \Mem_reg[55][4]  ( .D(n4050), .CLK(clk), .Q(\Mem[55][4] ) );
  DFFPOSX1 \Mem_reg[55][3]  ( .D(n4049), .CLK(clk), .Q(\Mem[55][3] ) );
  DFFPOSX1 \Mem_reg[55][2]  ( .D(n4048), .CLK(clk), .Q(\Mem[55][2] ) );
  DFFPOSX1 \Mem_reg[55][1]  ( .D(n4047), .CLK(clk), .Q(\Mem[55][1] ) );
  DFFPOSX1 \Mem_reg[55][0]  ( .D(n4046), .CLK(clk), .Q(\Mem[55][0] ) );
  DFFPOSX1 \Mem_reg[54][31]  ( .D(n4045), .CLK(clk), .Q(\Mem[54][31] ) );
  DFFPOSX1 \Mem_reg[54][30]  ( .D(n4044), .CLK(clk), .Q(\Mem[54][30] ) );
  DFFPOSX1 \Mem_reg[54][29]  ( .D(n4043), .CLK(clk), .Q(\Mem[54][29] ) );
  DFFPOSX1 \Mem_reg[54][28]  ( .D(n4042), .CLK(clk), .Q(\Mem[54][28] ) );
  DFFPOSX1 \Mem_reg[54][27]  ( .D(n4041), .CLK(clk), .Q(\Mem[54][27] ) );
  DFFPOSX1 \Mem_reg[54][26]  ( .D(n4040), .CLK(clk), .Q(\Mem[54][26] ) );
  DFFPOSX1 \Mem_reg[54][25]  ( .D(n4039), .CLK(clk), .Q(\Mem[54][25] ) );
  DFFPOSX1 \Mem_reg[54][24]  ( .D(n4038), .CLK(clk), .Q(\Mem[54][24] ) );
  DFFPOSX1 \Mem_reg[54][23]  ( .D(n4037), .CLK(clk), .Q(\Mem[54][23] ) );
  DFFPOSX1 \Mem_reg[54][22]  ( .D(n4036), .CLK(clk), .Q(\Mem[54][22] ) );
  DFFPOSX1 \Mem_reg[54][21]  ( .D(n4035), .CLK(clk), .Q(\Mem[54][21] ) );
  DFFPOSX1 \Mem_reg[54][20]  ( .D(n4034), .CLK(clk), .Q(\Mem[54][20] ) );
  DFFPOSX1 \Mem_reg[54][19]  ( .D(n4033), .CLK(clk), .Q(\Mem[54][19] ) );
  DFFPOSX1 \Mem_reg[54][18]  ( .D(n4032), .CLK(clk), .Q(\Mem[54][18] ) );
  DFFPOSX1 \Mem_reg[54][17]  ( .D(n4031), .CLK(clk), .Q(\Mem[54][17] ) );
  DFFPOSX1 \Mem_reg[54][16]  ( .D(n4030), .CLK(clk), .Q(\Mem[54][16] ) );
  DFFPOSX1 \Mem_reg[54][15]  ( .D(n4029), .CLK(clk), .Q(\Mem[54][15] ) );
  DFFPOSX1 \Mem_reg[54][14]  ( .D(n4028), .CLK(clk), .Q(\Mem[54][14] ) );
  DFFPOSX1 \Mem_reg[54][13]  ( .D(n4027), .CLK(clk), .Q(\Mem[54][13] ) );
  DFFPOSX1 \Mem_reg[54][12]  ( .D(n4026), .CLK(clk), .Q(\Mem[54][12] ) );
  DFFPOSX1 \Mem_reg[54][11]  ( .D(n4025), .CLK(clk), .Q(\Mem[54][11] ) );
  DFFPOSX1 \Mem_reg[54][10]  ( .D(n4024), .CLK(clk), .Q(\Mem[54][10] ) );
  DFFPOSX1 \Mem_reg[54][9]  ( .D(n4023), .CLK(clk), .Q(\Mem[54][9] ) );
  DFFPOSX1 \Mem_reg[54][8]  ( .D(n4022), .CLK(clk), .Q(\Mem[54][8] ) );
  DFFPOSX1 \Mem_reg[54][7]  ( .D(n4021), .CLK(clk), .Q(\Mem[54][7] ) );
  DFFPOSX1 \Mem_reg[54][6]  ( .D(n4020), .CLK(clk), .Q(\Mem[54][6] ) );
  DFFPOSX1 \Mem_reg[54][5]  ( .D(n4019), .CLK(clk), .Q(\Mem[54][5] ) );
  DFFPOSX1 \Mem_reg[54][4]  ( .D(n4018), .CLK(clk), .Q(\Mem[54][4] ) );
  DFFPOSX1 \Mem_reg[54][3]  ( .D(n4017), .CLK(clk), .Q(\Mem[54][3] ) );
  DFFPOSX1 \Mem_reg[54][2]  ( .D(n4016), .CLK(clk), .Q(\Mem[54][2] ) );
  DFFPOSX1 \Mem_reg[54][1]  ( .D(n4015), .CLK(clk), .Q(\Mem[54][1] ) );
  DFFPOSX1 \Mem_reg[54][0]  ( .D(n4014), .CLK(clk), .Q(\Mem[54][0] ) );
  DFFPOSX1 \Mem_reg[53][31]  ( .D(n4013), .CLK(clk), .Q(\Mem[53][31] ) );
  DFFPOSX1 \Mem_reg[53][30]  ( .D(n4012), .CLK(clk), .Q(\Mem[53][30] ) );
  DFFPOSX1 \Mem_reg[53][29]  ( .D(n4011), .CLK(clk), .Q(\Mem[53][29] ) );
  DFFPOSX1 \Mem_reg[53][28]  ( .D(n4010), .CLK(clk), .Q(\Mem[53][28] ) );
  DFFPOSX1 \Mem_reg[53][27]  ( .D(n4009), .CLK(clk), .Q(\Mem[53][27] ) );
  DFFPOSX1 \Mem_reg[53][26]  ( .D(n4008), .CLK(clk), .Q(\Mem[53][26] ) );
  DFFPOSX1 \Mem_reg[53][25]  ( .D(n4007), .CLK(clk), .Q(\Mem[53][25] ) );
  DFFPOSX1 \Mem_reg[53][24]  ( .D(n4006), .CLK(clk), .Q(\Mem[53][24] ) );
  DFFPOSX1 \Mem_reg[53][23]  ( .D(n4005), .CLK(clk), .Q(\Mem[53][23] ) );
  DFFPOSX1 \Mem_reg[53][22]  ( .D(n4004), .CLK(clk), .Q(\Mem[53][22] ) );
  DFFPOSX1 \Mem_reg[53][21]  ( .D(n4003), .CLK(clk), .Q(\Mem[53][21] ) );
  DFFPOSX1 \Mem_reg[53][20]  ( .D(n4002), .CLK(clk), .Q(\Mem[53][20] ) );
  DFFPOSX1 \Mem_reg[53][19]  ( .D(n4001), .CLK(clk), .Q(\Mem[53][19] ) );
  DFFPOSX1 \Mem_reg[53][18]  ( .D(n4000), .CLK(clk), .Q(\Mem[53][18] ) );
  DFFPOSX1 \Mem_reg[53][17]  ( .D(n3999), .CLK(clk), .Q(\Mem[53][17] ) );
  DFFPOSX1 \Mem_reg[53][16]  ( .D(n3998), .CLK(clk), .Q(\Mem[53][16] ) );
  DFFPOSX1 \Mem_reg[53][15]  ( .D(n3997), .CLK(clk), .Q(\Mem[53][15] ) );
  DFFPOSX1 \Mem_reg[53][14]  ( .D(n3996), .CLK(clk), .Q(\Mem[53][14] ) );
  DFFPOSX1 \Mem_reg[53][13]  ( .D(n3995), .CLK(clk), .Q(\Mem[53][13] ) );
  DFFPOSX1 \Mem_reg[53][12]  ( .D(n3994), .CLK(clk), .Q(\Mem[53][12] ) );
  DFFPOSX1 \Mem_reg[53][11]  ( .D(n3993), .CLK(clk), .Q(\Mem[53][11] ) );
  DFFPOSX1 \Mem_reg[53][10]  ( .D(n3992), .CLK(clk), .Q(\Mem[53][10] ) );
  DFFPOSX1 \Mem_reg[53][9]  ( .D(n3991), .CLK(clk), .Q(\Mem[53][9] ) );
  DFFPOSX1 \Mem_reg[53][8]  ( .D(n3990), .CLK(clk), .Q(\Mem[53][8] ) );
  DFFPOSX1 \Mem_reg[53][7]  ( .D(n3989), .CLK(clk), .Q(\Mem[53][7] ) );
  DFFPOSX1 \Mem_reg[53][6]  ( .D(n3988), .CLK(clk), .Q(\Mem[53][6] ) );
  DFFPOSX1 \Mem_reg[53][5]  ( .D(n3987), .CLK(clk), .Q(\Mem[53][5] ) );
  DFFPOSX1 \Mem_reg[53][4]  ( .D(n3986), .CLK(clk), .Q(\Mem[53][4] ) );
  DFFPOSX1 \Mem_reg[53][3]  ( .D(n3985), .CLK(clk), .Q(\Mem[53][3] ) );
  DFFPOSX1 \Mem_reg[53][2]  ( .D(n3984), .CLK(clk), .Q(\Mem[53][2] ) );
  DFFPOSX1 \Mem_reg[53][1]  ( .D(n3983), .CLK(clk), .Q(\Mem[53][1] ) );
  DFFPOSX1 \Mem_reg[53][0]  ( .D(n3982), .CLK(clk), .Q(\Mem[53][0] ) );
  DFFPOSX1 \Mem_reg[52][31]  ( .D(n3981), .CLK(clk), .Q(\Mem[52][31] ) );
  DFFPOSX1 \Mem_reg[52][30]  ( .D(n3980), .CLK(clk), .Q(\Mem[52][30] ) );
  DFFPOSX1 \Mem_reg[52][29]  ( .D(n3979), .CLK(clk), .Q(\Mem[52][29] ) );
  DFFPOSX1 \Mem_reg[52][28]  ( .D(n3978), .CLK(clk), .Q(\Mem[52][28] ) );
  DFFPOSX1 \Mem_reg[52][27]  ( .D(n3977), .CLK(clk), .Q(\Mem[52][27] ) );
  DFFPOSX1 \Mem_reg[52][26]  ( .D(n3976), .CLK(clk), .Q(\Mem[52][26] ) );
  DFFPOSX1 \Mem_reg[52][25]  ( .D(n3975), .CLK(clk), .Q(\Mem[52][25] ) );
  DFFPOSX1 \Mem_reg[52][24]  ( .D(n3974), .CLK(clk), .Q(\Mem[52][24] ) );
  DFFPOSX1 \Mem_reg[52][23]  ( .D(n3973), .CLK(clk), .Q(\Mem[52][23] ) );
  DFFPOSX1 \Mem_reg[52][22]  ( .D(n3972), .CLK(clk), .Q(\Mem[52][22] ) );
  DFFPOSX1 \Mem_reg[52][21]  ( .D(n3971), .CLK(clk), .Q(\Mem[52][21] ) );
  DFFPOSX1 \Mem_reg[52][20]  ( .D(n3970), .CLK(clk), .Q(\Mem[52][20] ) );
  DFFPOSX1 \Mem_reg[52][19]  ( .D(n3969), .CLK(clk), .Q(\Mem[52][19] ) );
  DFFPOSX1 \Mem_reg[52][18]  ( .D(n3968), .CLK(clk), .Q(\Mem[52][18] ) );
  DFFPOSX1 \Mem_reg[52][17]  ( .D(n3967), .CLK(clk), .Q(\Mem[52][17] ) );
  DFFPOSX1 \Mem_reg[52][16]  ( .D(n3966), .CLK(clk), .Q(\Mem[52][16] ) );
  DFFPOSX1 \Mem_reg[52][15]  ( .D(n3965), .CLK(clk), .Q(\Mem[52][15] ) );
  DFFPOSX1 \Mem_reg[52][14]  ( .D(n3964), .CLK(clk), .Q(\Mem[52][14] ) );
  DFFPOSX1 \Mem_reg[52][13]  ( .D(n3963), .CLK(clk), .Q(\Mem[52][13] ) );
  DFFPOSX1 \Mem_reg[52][12]  ( .D(n3962), .CLK(clk), .Q(\Mem[52][12] ) );
  DFFPOSX1 \Mem_reg[52][11]  ( .D(n3961), .CLK(clk), .Q(\Mem[52][11] ) );
  DFFPOSX1 \Mem_reg[52][10]  ( .D(n3960), .CLK(clk), .Q(\Mem[52][10] ) );
  DFFPOSX1 \Mem_reg[52][9]  ( .D(n3959), .CLK(clk), .Q(\Mem[52][9] ) );
  DFFPOSX1 \Mem_reg[52][8]  ( .D(n3958), .CLK(clk), .Q(\Mem[52][8] ) );
  DFFPOSX1 \Mem_reg[52][7]  ( .D(n3957), .CLK(clk), .Q(\Mem[52][7] ) );
  DFFPOSX1 \Mem_reg[52][6]  ( .D(n3956), .CLK(clk), .Q(\Mem[52][6] ) );
  DFFPOSX1 \Mem_reg[52][5]  ( .D(n3955), .CLK(clk), .Q(\Mem[52][5] ) );
  DFFPOSX1 \Mem_reg[52][4]  ( .D(n3954), .CLK(clk), .Q(\Mem[52][4] ) );
  DFFPOSX1 \Mem_reg[52][3]  ( .D(n3953), .CLK(clk), .Q(\Mem[52][3] ) );
  DFFPOSX1 \Mem_reg[52][2]  ( .D(n3952), .CLK(clk), .Q(\Mem[52][2] ) );
  DFFPOSX1 \Mem_reg[52][1]  ( .D(n3951), .CLK(clk), .Q(\Mem[52][1] ) );
  DFFPOSX1 \Mem_reg[52][0]  ( .D(n3950), .CLK(clk), .Q(\Mem[52][0] ) );
  DFFPOSX1 \Mem_reg[51][31]  ( .D(n3949), .CLK(clk), .Q(\Mem[51][31] ) );
  DFFPOSX1 \Mem_reg[51][30]  ( .D(n3948), .CLK(clk), .Q(\Mem[51][30] ) );
  DFFPOSX1 \Mem_reg[51][29]  ( .D(n3947), .CLK(clk), .Q(\Mem[51][29] ) );
  DFFPOSX1 \Mem_reg[51][28]  ( .D(n3946), .CLK(clk), .Q(\Mem[51][28] ) );
  DFFPOSX1 \Mem_reg[51][27]  ( .D(n3945), .CLK(clk), .Q(\Mem[51][27] ) );
  DFFPOSX1 \Mem_reg[51][26]  ( .D(n3944), .CLK(clk), .Q(\Mem[51][26] ) );
  DFFPOSX1 \Mem_reg[51][25]  ( .D(n3943), .CLK(clk), .Q(\Mem[51][25] ) );
  DFFPOSX1 \Mem_reg[51][24]  ( .D(n3942), .CLK(clk), .Q(\Mem[51][24] ) );
  DFFPOSX1 \Mem_reg[51][23]  ( .D(n3941), .CLK(clk), .Q(\Mem[51][23] ) );
  DFFPOSX1 \Mem_reg[51][22]  ( .D(n3940), .CLK(clk), .Q(\Mem[51][22] ) );
  DFFPOSX1 \Mem_reg[51][21]  ( .D(n3939), .CLK(clk), .Q(\Mem[51][21] ) );
  DFFPOSX1 \Mem_reg[51][20]  ( .D(n3938), .CLK(clk), .Q(\Mem[51][20] ) );
  DFFPOSX1 \Mem_reg[51][19]  ( .D(n3937), .CLK(clk), .Q(\Mem[51][19] ) );
  DFFPOSX1 \Mem_reg[51][18]  ( .D(n3936), .CLK(clk), .Q(\Mem[51][18] ) );
  DFFPOSX1 \Mem_reg[51][17]  ( .D(n3935), .CLK(clk), .Q(\Mem[51][17] ) );
  DFFPOSX1 \Mem_reg[51][16]  ( .D(n3934), .CLK(clk), .Q(\Mem[51][16] ) );
  DFFPOSX1 \Mem_reg[51][15]  ( .D(n3933), .CLK(clk), .Q(\Mem[51][15] ) );
  DFFPOSX1 \Mem_reg[51][14]  ( .D(n3932), .CLK(clk), .Q(\Mem[51][14] ) );
  DFFPOSX1 \Mem_reg[51][13]  ( .D(n3931), .CLK(clk), .Q(\Mem[51][13] ) );
  DFFPOSX1 \Mem_reg[51][12]  ( .D(n3930), .CLK(clk), .Q(\Mem[51][12] ) );
  DFFPOSX1 \Mem_reg[51][11]  ( .D(n3929), .CLK(clk), .Q(\Mem[51][11] ) );
  DFFPOSX1 \Mem_reg[51][10]  ( .D(n3928), .CLK(clk), .Q(\Mem[51][10] ) );
  DFFPOSX1 \Mem_reg[51][9]  ( .D(n3927), .CLK(clk), .Q(\Mem[51][9] ) );
  DFFPOSX1 \Mem_reg[51][8]  ( .D(n3926), .CLK(clk), .Q(\Mem[51][8] ) );
  DFFPOSX1 \Mem_reg[51][7]  ( .D(n3925), .CLK(clk), .Q(\Mem[51][7] ) );
  DFFPOSX1 \Mem_reg[51][6]  ( .D(n3924), .CLK(clk), .Q(\Mem[51][6] ) );
  DFFPOSX1 \Mem_reg[51][5]  ( .D(n3923), .CLK(clk), .Q(\Mem[51][5] ) );
  DFFPOSX1 \Mem_reg[51][4]  ( .D(n3922), .CLK(clk), .Q(\Mem[51][4] ) );
  DFFPOSX1 \Mem_reg[51][3]  ( .D(n3921), .CLK(clk), .Q(\Mem[51][3] ) );
  DFFPOSX1 \Mem_reg[51][2]  ( .D(n3920), .CLK(clk), .Q(\Mem[51][2] ) );
  DFFPOSX1 \Mem_reg[51][1]  ( .D(n3919), .CLK(clk), .Q(\Mem[51][1] ) );
  DFFPOSX1 \Mem_reg[51][0]  ( .D(n3918), .CLK(clk), .Q(\Mem[51][0] ) );
  DFFPOSX1 \Mem_reg[50][31]  ( .D(n3917), .CLK(clk), .Q(\Mem[50][31] ) );
  DFFPOSX1 \Mem_reg[50][30]  ( .D(n3916), .CLK(clk), .Q(\Mem[50][30] ) );
  DFFPOSX1 \Mem_reg[50][29]  ( .D(n3915), .CLK(clk), .Q(\Mem[50][29] ) );
  DFFPOSX1 \Mem_reg[50][28]  ( .D(n3914), .CLK(clk), .Q(\Mem[50][28] ) );
  DFFPOSX1 \Mem_reg[50][27]  ( .D(n3913), .CLK(clk), .Q(\Mem[50][27] ) );
  DFFPOSX1 \Mem_reg[50][26]  ( .D(n3912), .CLK(clk), .Q(\Mem[50][26] ) );
  DFFPOSX1 \Mem_reg[50][25]  ( .D(n3911), .CLK(clk), .Q(\Mem[50][25] ) );
  DFFPOSX1 \Mem_reg[50][24]  ( .D(n3910), .CLK(clk), .Q(\Mem[50][24] ) );
  DFFPOSX1 \Mem_reg[50][23]  ( .D(n3909), .CLK(clk), .Q(\Mem[50][23] ) );
  DFFPOSX1 \Mem_reg[50][22]  ( .D(n3908), .CLK(clk), .Q(\Mem[50][22] ) );
  DFFPOSX1 \Mem_reg[50][21]  ( .D(n3907), .CLK(clk), .Q(\Mem[50][21] ) );
  DFFPOSX1 \Mem_reg[50][20]  ( .D(n3906), .CLK(clk), .Q(\Mem[50][20] ) );
  DFFPOSX1 \Mem_reg[50][19]  ( .D(n3905), .CLK(clk), .Q(\Mem[50][19] ) );
  DFFPOSX1 \Mem_reg[50][18]  ( .D(n3904), .CLK(clk), .Q(\Mem[50][18] ) );
  DFFPOSX1 \Mem_reg[50][17]  ( .D(n3903), .CLK(clk), .Q(\Mem[50][17] ) );
  DFFPOSX1 \Mem_reg[50][16]  ( .D(n3902), .CLK(clk), .Q(\Mem[50][16] ) );
  DFFPOSX1 \Mem_reg[50][15]  ( .D(n3901), .CLK(clk), .Q(\Mem[50][15] ) );
  DFFPOSX1 \Mem_reg[50][14]  ( .D(n3900), .CLK(clk), .Q(\Mem[50][14] ) );
  DFFPOSX1 \Mem_reg[50][13]  ( .D(n3899), .CLK(clk), .Q(\Mem[50][13] ) );
  DFFPOSX1 \Mem_reg[50][12]  ( .D(n3898), .CLK(clk), .Q(\Mem[50][12] ) );
  DFFPOSX1 \Mem_reg[50][11]  ( .D(n3897), .CLK(clk), .Q(\Mem[50][11] ) );
  DFFPOSX1 \Mem_reg[50][10]  ( .D(n3896), .CLK(clk), .Q(\Mem[50][10] ) );
  DFFPOSX1 \Mem_reg[50][9]  ( .D(n3895), .CLK(clk), .Q(\Mem[50][9] ) );
  DFFPOSX1 \Mem_reg[50][8]  ( .D(n3894), .CLK(clk), .Q(\Mem[50][8] ) );
  DFFPOSX1 \Mem_reg[50][7]  ( .D(n3893), .CLK(clk), .Q(\Mem[50][7] ) );
  DFFPOSX1 \Mem_reg[50][6]  ( .D(n3892), .CLK(clk), .Q(\Mem[50][6] ) );
  DFFPOSX1 \Mem_reg[50][5]  ( .D(n3891), .CLK(clk), .Q(\Mem[50][5] ) );
  DFFPOSX1 \Mem_reg[50][4]  ( .D(n3890), .CLK(clk), .Q(\Mem[50][4] ) );
  DFFPOSX1 \Mem_reg[50][3]  ( .D(n3889), .CLK(clk), .Q(\Mem[50][3] ) );
  DFFPOSX1 \Mem_reg[50][2]  ( .D(n3888), .CLK(clk), .Q(\Mem[50][2] ) );
  DFFPOSX1 \Mem_reg[50][1]  ( .D(n3887), .CLK(clk), .Q(\Mem[50][1] ) );
  DFFPOSX1 \Mem_reg[50][0]  ( .D(n3886), .CLK(clk), .Q(\Mem[50][0] ) );
  DFFPOSX1 \Mem_reg[49][31]  ( .D(n3885), .CLK(clk), .Q(\Mem[49][31] ) );
  DFFPOSX1 \Mem_reg[49][30]  ( .D(n3884), .CLK(clk), .Q(\Mem[49][30] ) );
  DFFPOSX1 \Mem_reg[49][29]  ( .D(n3883), .CLK(clk), .Q(\Mem[49][29] ) );
  DFFPOSX1 \Mem_reg[49][28]  ( .D(n3882), .CLK(clk), .Q(\Mem[49][28] ) );
  DFFPOSX1 \Mem_reg[49][27]  ( .D(n3881), .CLK(clk), .Q(\Mem[49][27] ) );
  DFFPOSX1 \Mem_reg[49][26]  ( .D(n3880), .CLK(clk), .Q(\Mem[49][26] ) );
  DFFPOSX1 \Mem_reg[49][25]  ( .D(n3879), .CLK(clk), .Q(\Mem[49][25] ) );
  DFFPOSX1 \Mem_reg[49][24]  ( .D(n3878), .CLK(clk), .Q(\Mem[49][24] ) );
  DFFPOSX1 \Mem_reg[49][23]  ( .D(n3877), .CLK(clk), .Q(\Mem[49][23] ) );
  DFFPOSX1 \Mem_reg[49][22]  ( .D(n3876), .CLK(clk), .Q(\Mem[49][22] ) );
  DFFPOSX1 \Mem_reg[49][21]  ( .D(n3875), .CLK(clk), .Q(\Mem[49][21] ) );
  DFFPOSX1 \Mem_reg[49][20]  ( .D(n3874), .CLK(clk), .Q(\Mem[49][20] ) );
  DFFPOSX1 \Mem_reg[49][19]  ( .D(n3873), .CLK(clk), .Q(\Mem[49][19] ) );
  DFFPOSX1 \Mem_reg[49][18]  ( .D(n3872), .CLK(clk), .Q(\Mem[49][18] ) );
  DFFPOSX1 \Mem_reg[49][17]  ( .D(n3871), .CLK(clk), .Q(\Mem[49][17] ) );
  DFFPOSX1 \Mem_reg[49][16]  ( .D(n3870), .CLK(clk), .Q(\Mem[49][16] ) );
  DFFPOSX1 \Mem_reg[49][15]  ( .D(n3869), .CLK(clk), .Q(\Mem[49][15] ) );
  DFFPOSX1 \Mem_reg[49][14]  ( .D(n3868), .CLK(clk), .Q(\Mem[49][14] ) );
  DFFPOSX1 \Mem_reg[49][13]  ( .D(n3867), .CLK(clk), .Q(\Mem[49][13] ) );
  DFFPOSX1 \Mem_reg[49][12]  ( .D(n3866), .CLK(clk), .Q(\Mem[49][12] ) );
  DFFPOSX1 \Mem_reg[49][11]  ( .D(n3865), .CLK(clk), .Q(\Mem[49][11] ) );
  DFFPOSX1 \Mem_reg[49][10]  ( .D(n3864), .CLK(clk), .Q(\Mem[49][10] ) );
  DFFPOSX1 \Mem_reg[49][9]  ( .D(n3863), .CLK(clk), .Q(\Mem[49][9] ) );
  DFFPOSX1 \Mem_reg[49][8]  ( .D(n3862), .CLK(clk), .Q(\Mem[49][8] ) );
  DFFPOSX1 \Mem_reg[49][7]  ( .D(n3861), .CLK(clk), .Q(\Mem[49][7] ) );
  DFFPOSX1 \Mem_reg[49][6]  ( .D(n3860), .CLK(clk), .Q(\Mem[49][6] ) );
  DFFPOSX1 \Mem_reg[49][5]  ( .D(n3859), .CLK(clk), .Q(\Mem[49][5] ) );
  DFFPOSX1 \Mem_reg[49][4]  ( .D(n3858), .CLK(clk), .Q(\Mem[49][4] ) );
  DFFPOSX1 \Mem_reg[49][3]  ( .D(n3857), .CLK(clk), .Q(\Mem[49][3] ) );
  DFFPOSX1 \Mem_reg[49][2]  ( .D(n3856), .CLK(clk), .Q(\Mem[49][2] ) );
  DFFPOSX1 \Mem_reg[49][1]  ( .D(n3855), .CLK(clk), .Q(\Mem[49][1] ) );
  DFFPOSX1 \Mem_reg[49][0]  ( .D(n3854), .CLK(clk), .Q(\Mem[49][0] ) );
  DFFPOSX1 \Mem_reg[48][31]  ( .D(n3853), .CLK(clk), .Q(\Mem[48][31] ) );
  DFFPOSX1 \Mem_reg[48][30]  ( .D(n3852), .CLK(clk), .Q(\Mem[48][30] ) );
  DFFPOSX1 \Mem_reg[48][29]  ( .D(n3851), .CLK(clk), .Q(\Mem[48][29] ) );
  DFFPOSX1 \Mem_reg[48][28]  ( .D(n3850), .CLK(clk), .Q(\Mem[48][28] ) );
  DFFPOSX1 \Mem_reg[48][27]  ( .D(n3849), .CLK(clk), .Q(\Mem[48][27] ) );
  DFFPOSX1 \Mem_reg[48][26]  ( .D(n3848), .CLK(clk), .Q(\Mem[48][26] ) );
  DFFPOSX1 \Mem_reg[48][25]  ( .D(n3847), .CLK(clk), .Q(\Mem[48][25] ) );
  DFFPOSX1 \Mem_reg[48][24]  ( .D(n3846), .CLK(clk), .Q(\Mem[48][24] ) );
  DFFPOSX1 \Mem_reg[48][23]  ( .D(n3845), .CLK(clk), .Q(\Mem[48][23] ) );
  DFFPOSX1 \Mem_reg[48][22]  ( .D(n3844), .CLK(clk), .Q(\Mem[48][22] ) );
  DFFPOSX1 \Mem_reg[48][21]  ( .D(n3843), .CLK(clk), .Q(\Mem[48][21] ) );
  DFFPOSX1 \Mem_reg[48][20]  ( .D(n3842), .CLK(clk), .Q(\Mem[48][20] ) );
  DFFPOSX1 \Mem_reg[48][19]  ( .D(n3841), .CLK(clk), .Q(\Mem[48][19] ) );
  DFFPOSX1 \Mem_reg[48][18]  ( .D(n3840), .CLK(clk), .Q(\Mem[48][18] ) );
  DFFPOSX1 \Mem_reg[48][17]  ( .D(n3839), .CLK(clk), .Q(\Mem[48][17] ) );
  DFFPOSX1 \Mem_reg[48][16]  ( .D(n3838), .CLK(clk), .Q(\Mem[48][16] ) );
  DFFPOSX1 \Mem_reg[48][15]  ( .D(n3837), .CLK(clk), .Q(\Mem[48][15] ) );
  DFFPOSX1 \Mem_reg[48][14]  ( .D(n3836), .CLK(clk), .Q(\Mem[48][14] ) );
  DFFPOSX1 \Mem_reg[48][13]  ( .D(n3835), .CLK(clk), .Q(\Mem[48][13] ) );
  DFFPOSX1 \Mem_reg[48][12]  ( .D(n3834), .CLK(clk), .Q(\Mem[48][12] ) );
  DFFPOSX1 \Mem_reg[48][11]  ( .D(n3833), .CLK(clk), .Q(\Mem[48][11] ) );
  DFFPOSX1 \Mem_reg[48][10]  ( .D(n3832), .CLK(clk), .Q(\Mem[48][10] ) );
  DFFPOSX1 \Mem_reg[48][9]  ( .D(n3831), .CLK(clk), .Q(\Mem[48][9] ) );
  DFFPOSX1 \Mem_reg[48][8]  ( .D(n3830), .CLK(clk), .Q(\Mem[48][8] ) );
  DFFPOSX1 \Mem_reg[48][7]  ( .D(n3829), .CLK(clk), .Q(\Mem[48][7] ) );
  DFFPOSX1 \Mem_reg[48][6]  ( .D(n3828), .CLK(clk), .Q(\Mem[48][6] ) );
  DFFPOSX1 \Mem_reg[48][5]  ( .D(n3827), .CLK(clk), .Q(\Mem[48][5] ) );
  DFFPOSX1 \Mem_reg[48][4]  ( .D(n3826), .CLK(clk), .Q(\Mem[48][4] ) );
  DFFPOSX1 \Mem_reg[48][3]  ( .D(n3825), .CLK(clk), .Q(\Mem[48][3] ) );
  DFFPOSX1 \Mem_reg[48][2]  ( .D(n3824), .CLK(clk), .Q(\Mem[48][2] ) );
  DFFPOSX1 \Mem_reg[48][1]  ( .D(n3823), .CLK(clk), .Q(\Mem[48][1] ) );
  DFFPOSX1 \Mem_reg[48][0]  ( .D(n3822), .CLK(clk), .Q(\Mem[48][0] ) );
  DFFPOSX1 \Mem_reg[47][31]  ( .D(n3821), .CLK(clk), .Q(\Mem[47][31] ) );
  DFFPOSX1 \Mem_reg[47][30]  ( .D(n3820), .CLK(clk), .Q(\Mem[47][30] ) );
  DFFPOSX1 \Mem_reg[47][29]  ( .D(n3819), .CLK(clk), .Q(\Mem[47][29] ) );
  DFFPOSX1 \Mem_reg[47][28]  ( .D(n3818), .CLK(clk), .Q(\Mem[47][28] ) );
  DFFPOSX1 \Mem_reg[47][27]  ( .D(n3817), .CLK(clk), .Q(\Mem[47][27] ) );
  DFFPOSX1 \Mem_reg[47][26]  ( .D(n3816), .CLK(clk), .Q(\Mem[47][26] ) );
  DFFPOSX1 \Mem_reg[47][25]  ( .D(n3815), .CLK(clk), .Q(\Mem[47][25] ) );
  DFFPOSX1 \Mem_reg[47][24]  ( .D(n3814), .CLK(clk), .Q(\Mem[47][24] ) );
  DFFPOSX1 \Mem_reg[47][23]  ( .D(n3813), .CLK(clk), .Q(\Mem[47][23] ) );
  DFFPOSX1 \Mem_reg[47][22]  ( .D(n3812), .CLK(clk), .Q(\Mem[47][22] ) );
  DFFPOSX1 \Mem_reg[47][21]  ( .D(n3811), .CLK(clk), .Q(\Mem[47][21] ) );
  DFFPOSX1 \Mem_reg[47][20]  ( .D(n3810), .CLK(clk), .Q(\Mem[47][20] ) );
  DFFPOSX1 \Mem_reg[47][19]  ( .D(n3809), .CLK(clk), .Q(\Mem[47][19] ) );
  DFFPOSX1 \Mem_reg[47][18]  ( .D(n3808), .CLK(clk), .Q(\Mem[47][18] ) );
  DFFPOSX1 \Mem_reg[47][17]  ( .D(n3807), .CLK(clk), .Q(\Mem[47][17] ) );
  DFFPOSX1 \Mem_reg[47][16]  ( .D(n3806), .CLK(clk), .Q(\Mem[47][16] ) );
  DFFPOSX1 \Mem_reg[47][15]  ( .D(n3805), .CLK(clk), .Q(\Mem[47][15] ) );
  DFFPOSX1 \Mem_reg[47][14]  ( .D(n3804), .CLK(clk), .Q(\Mem[47][14] ) );
  DFFPOSX1 \Mem_reg[47][13]  ( .D(n3803), .CLK(clk), .Q(\Mem[47][13] ) );
  DFFPOSX1 \Mem_reg[47][12]  ( .D(n3802), .CLK(clk), .Q(\Mem[47][12] ) );
  DFFPOSX1 \Mem_reg[47][11]  ( .D(n3801), .CLK(clk), .Q(\Mem[47][11] ) );
  DFFPOSX1 \Mem_reg[47][10]  ( .D(n3800), .CLK(clk), .Q(\Mem[47][10] ) );
  DFFPOSX1 \Mem_reg[47][9]  ( .D(n3799), .CLK(clk), .Q(\Mem[47][9] ) );
  DFFPOSX1 \Mem_reg[47][8]  ( .D(n3798), .CLK(clk), .Q(\Mem[47][8] ) );
  DFFPOSX1 \Mem_reg[47][7]  ( .D(n3797), .CLK(clk), .Q(\Mem[47][7] ) );
  DFFPOSX1 \Mem_reg[47][6]  ( .D(n3796), .CLK(clk), .Q(\Mem[47][6] ) );
  DFFPOSX1 \Mem_reg[47][5]  ( .D(n3795), .CLK(clk), .Q(\Mem[47][5] ) );
  DFFPOSX1 \Mem_reg[47][4]  ( .D(n3794), .CLK(clk), .Q(\Mem[47][4] ) );
  DFFPOSX1 \Mem_reg[47][3]  ( .D(n3793), .CLK(clk), .Q(\Mem[47][3] ) );
  DFFPOSX1 \Mem_reg[47][2]  ( .D(n3792), .CLK(clk), .Q(\Mem[47][2] ) );
  DFFPOSX1 \Mem_reg[47][1]  ( .D(n3791), .CLK(clk), .Q(\Mem[47][1] ) );
  DFFPOSX1 \Mem_reg[47][0]  ( .D(n3790), .CLK(clk), .Q(\Mem[47][0] ) );
  DFFPOSX1 \Mem_reg[46][31]  ( .D(n3789), .CLK(clk), .Q(\Mem[46][31] ) );
  DFFPOSX1 \Mem_reg[46][30]  ( .D(n3788), .CLK(clk), .Q(\Mem[46][30] ) );
  DFFPOSX1 \Mem_reg[46][29]  ( .D(n3787), .CLK(clk), .Q(\Mem[46][29] ) );
  DFFPOSX1 \Mem_reg[46][28]  ( .D(n3786), .CLK(clk), .Q(\Mem[46][28] ) );
  DFFPOSX1 \Mem_reg[46][27]  ( .D(n3785), .CLK(clk), .Q(\Mem[46][27] ) );
  DFFPOSX1 \Mem_reg[46][26]  ( .D(n3784), .CLK(clk), .Q(\Mem[46][26] ) );
  DFFPOSX1 \Mem_reg[46][25]  ( .D(n3783), .CLK(clk), .Q(\Mem[46][25] ) );
  DFFPOSX1 \Mem_reg[46][24]  ( .D(n3782), .CLK(clk), .Q(\Mem[46][24] ) );
  DFFPOSX1 \Mem_reg[46][23]  ( .D(n3781), .CLK(clk), .Q(\Mem[46][23] ) );
  DFFPOSX1 \Mem_reg[46][22]  ( .D(n3780), .CLK(clk), .Q(\Mem[46][22] ) );
  DFFPOSX1 \Mem_reg[46][21]  ( .D(n3779), .CLK(clk), .Q(\Mem[46][21] ) );
  DFFPOSX1 \Mem_reg[46][20]  ( .D(n3778), .CLK(clk), .Q(\Mem[46][20] ) );
  DFFPOSX1 \Mem_reg[46][19]  ( .D(n3777), .CLK(clk), .Q(\Mem[46][19] ) );
  DFFPOSX1 \Mem_reg[46][18]  ( .D(n3776), .CLK(clk), .Q(\Mem[46][18] ) );
  DFFPOSX1 \Mem_reg[46][17]  ( .D(n3775), .CLK(clk), .Q(\Mem[46][17] ) );
  DFFPOSX1 \Mem_reg[46][16]  ( .D(n3774), .CLK(clk), .Q(\Mem[46][16] ) );
  DFFPOSX1 \Mem_reg[46][15]  ( .D(n3773), .CLK(clk), .Q(\Mem[46][15] ) );
  DFFPOSX1 \Mem_reg[46][14]  ( .D(n3772), .CLK(clk), .Q(\Mem[46][14] ) );
  DFFPOSX1 \Mem_reg[46][13]  ( .D(n3771), .CLK(clk), .Q(\Mem[46][13] ) );
  DFFPOSX1 \Mem_reg[46][12]  ( .D(n3770), .CLK(clk), .Q(\Mem[46][12] ) );
  DFFPOSX1 \Mem_reg[46][11]  ( .D(n3769), .CLK(clk), .Q(\Mem[46][11] ) );
  DFFPOSX1 \Mem_reg[46][10]  ( .D(n3768), .CLK(clk), .Q(\Mem[46][10] ) );
  DFFPOSX1 \Mem_reg[46][9]  ( .D(n3767), .CLK(clk), .Q(\Mem[46][9] ) );
  DFFPOSX1 \Mem_reg[46][8]  ( .D(n3766), .CLK(clk), .Q(\Mem[46][8] ) );
  DFFPOSX1 \Mem_reg[46][7]  ( .D(n3765), .CLK(clk), .Q(\Mem[46][7] ) );
  DFFPOSX1 \Mem_reg[46][6]  ( .D(n3764), .CLK(clk), .Q(\Mem[46][6] ) );
  DFFPOSX1 \Mem_reg[46][5]  ( .D(n3763), .CLK(clk), .Q(\Mem[46][5] ) );
  DFFPOSX1 \Mem_reg[46][4]  ( .D(n3762), .CLK(clk), .Q(\Mem[46][4] ) );
  DFFPOSX1 \Mem_reg[46][3]  ( .D(n3761), .CLK(clk), .Q(\Mem[46][3] ) );
  DFFPOSX1 \Mem_reg[46][2]  ( .D(n3760), .CLK(clk), .Q(\Mem[46][2] ) );
  DFFPOSX1 \Mem_reg[46][1]  ( .D(n3759), .CLK(clk), .Q(\Mem[46][1] ) );
  DFFPOSX1 \Mem_reg[46][0]  ( .D(n3758), .CLK(clk), .Q(\Mem[46][0] ) );
  DFFPOSX1 \Mem_reg[45][31]  ( .D(n3757), .CLK(clk), .Q(\Mem[45][31] ) );
  DFFPOSX1 \Mem_reg[45][30]  ( .D(n3756), .CLK(clk), .Q(\Mem[45][30] ) );
  DFFPOSX1 \Mem_reg[45][29]  ( .D(n3755), .CLK(clk), .Q(\Mem[45][29] ) );
  DFFPOSX1 \Mem_reg[45][28]  ( .D(n3754), .CLK(clk), .Q(\Mem[45][28] ) );
  DFFPOSX1 \Mem_reg[45][27]  ( .D(n3753), .CLK(clk), .Q(\Mem[45][27] ) );
  DFFPOSX1 \Mem_reg[45][26]  ( .D(n3752), .CLK(clk), .Q(\Mem[45][26] ) );
  DFFPOSX1 \Mem_reg[45][25]  ( .D(n3751), .CLK(clk), .Q(\Mem[45][25] ) );
  DFFPOSX1 \Mem_reg[45][24]  ( .D(n3750), .CLK(clk), .Q(\Mem[45][24] ) );
  DFFPOSX1 \Mem_reg[45][23]  ( .D(n3749), .CLK(clk), .Q(\Mem[45][23] ) );
  DFFPOSX1 \Mem_reg[45][22]  ( .D(n3748), .CLK(clk), .Q(\Mem[45][22] ) );
  DFFPOSX1 \Mem_reg[45][21]  ( .D(n3747), .CLK(clk), .Q(\Mem[45][21] ) );
  DFFPOSX1 \Mem_reg[45][20]  ( .D(n3746), .CLK(clk), .Q(\Mem[45][20] ) );
  DFFPOSX1 \Mem_reg[45][19]  ( .D(n3745), .CLK(clk), .Q(\Mem[45][19] ) );
  DFFPOSX1 \Mem_reg[45][18]  ( .D(n3744), .CLK(clk), .Q(\Mem[45][18] ) );
  DFFPOSX1 \Mem_reg[45][17]  ( .D(n3743), .CLK(clk), .Q(\Mem[45][17] ) );
  DFFPOSX1 \Mem_reg[45][16]  ( .D(n3742), .CLK(clk), .Q(\Mem[45][16] ) );
  DFFPOSX1 \Mem_reg[45][15]  ( .D(n3741), .CLK(clk), .Q(\Mem[45][15] ) );
  DFFPOSX1 \Mem_reg[45][14]  ( .D(n3740), .CLK(clk), .Q(\Mem[45][14] ) );
  DFFPOSX1 \Mem_reg[45][13]  ( .D(n3739), .CLK(clk), .Q(\Mem[45][13] ) );
  DFFPOSX1 \Mem_reg[45][12]  ( .D(n3738), .CLK(clk), .Q(\Mem[45][12] ) );
  DFFPOSX1 \Mem_reg[45][11]  ( .D(n3737), .CLK(clk), .Q(\Mem[45][11] ) );
  DFFPOSX1 \Mem_reg[45][10]  ( .D(n3736), .CLK(clk), .Q(\Mem[45][10] ) );
  DFFPOSX1 \Mem_reg[45][9]  ( .D(n3735), .CLK(clk), .Q(\Mem[45][9] ) );
  DFFPOSX1 \Mem_reg[45][8]  ( .D(n3734), .CLK(clk), .Q(\Mem[45][8] ) );
  DFFPOSX1 \Mem_reg[45][7]  ( .D(n3733), .CLK(clk), .Q(\Mem[45][7] ) );
  DFFPOSX1 \Mem_reg[45][6]  ( .D(n3732), .CLK(clk), .Q(\Mem[45][6] ) );
  DFFPOSX1 \Mem_reg[45][5]  ( .D(n3731), .CLK(clk), .Q(\Mem[45][5] ) );
  DFFPOSX1 \Mem_reg[45][4]  ( .D(n3730), .CLK(clk), .Q(\Mem[45][4] ) );
  DFFPOSX1 \Mem_reg[45][3]  ( .D(n3729), .CLK(clk), .Q(\Mem[45][3] ) );
  DFFPOSX1 \Mem_reg[45][2]  ( .D(n3728), .CLK(clk), .Q(\Mem[45][2] ) );
  DFFPOSX1 \Mem_reg[45][1]  ( .D(n3727), .CLK(clk), .Q(\Mem[45][1] ) );
  DFFPOSX1 \Mem_reg[45][0]  ( .D(n3726), .CLK(clk), .Q(\Mem[45][0] ) );
  DFFPOSX1 \Mem_reg[44][31]  ( .D(n3725), .CLK(clk), .Q(\Mem[44][31] ) );
  DFFPOSX1 \Mem_reg[44][30]  ( .D(n3724), .CLK(clk), .Q(\Mem[44][30] ) );
  DFFPOSX1 \Mem_reg[44][29]  ( .D(n3723), .CLK(clk), .Q(\Mem[44][29] ) );
  DFFPOSX1 \Mem_reg[44][28]  ( .D(n3722), .CLK(clk), .Q(\Mem[44][28] ) );
  DFFPOSX1 \Mem_reg[44][27]  ( .D(n3721), .CLK(clk), .Q(\Mem[44][27] ) );
  DFFPOSX1 \Mem_reg[44][26]  ( .D(n3720), .CLK(clk), .Q(\Mem[44][26] ) );
  DFFPOSX1 \Mem_reg[44][25]  ( .D(n3719), .CLK(clk), .Q(\Mem[44][25] ) );
  DFFPOSX1 \Mem_reg[44][24]  ( .D(n3718), .CLK(clk), .Q(\Mem[44][24] ) );
  DFFPOSX1 \Mem_reg[44][23]  ( .D(n3717), .CLK(clk), .Q(\Mem[44][23] ) );
  DFFPOSX1 \Mem_reg[44][22]  ( .D(n3716), .CLK(clk), .Q(\Mem[44][22] ) );
  DFFPOSX1 \Mem_reg[44][21]  ( .D(n3715), .CLK(clk), .Q(\Mem[44][21] ) );
  DFFPOSX1 \Mem_reg[44][20]  ( .D(n3714), .CLK(clk), .Q(\Mem[44][20] ) );
  DFFPOSX1 \Mem_reg[44][19]  ( .D(n3713), .CLK(clk), .Q(\Mem[44][19] ) );
  DFFPOSX1 \Mem_reg[44][18]  ( .D(n3712), .CLK(clk), .Q(\Mem[44][18] ) );
  DFFPOSX1 \Mem_reg[44][17]  ( .D(n3711), .CLK(clk), .Q(\Mem[44][17] ) );
  DFFPOSX1 \Mem_reg[44][16]  ( .D(n3710), .CLK(clk), .Q(\Mem[44][16] ) );
  DFFPOSX1 \Mem_reg[44][15]  ( .D(n3709), .CLK(clk), .Q(\Mem[44][15] ) );
  DFFPOSX1 \Mem_reg[44][14]  ( .D(n3708), .CLK(clk), .Q(\Mem[44][14] ) );
  DFFPOSX1 \Mem_reg[44][13]  ( .D(n3707), .CLK(clk), .Q(\Mem[44][13] ) );
  DFFPOSX1 \Mem_reg[44][12]  ( .D(n3706), .CLK(clk), .Q(\Mem[44][12] ) );
  DFFPOSX1 \Mem_reg[44][11]  ( .D(n3705), .CLK(clk), .Q(\Mem[44][11] ) );
  DFFPOSX1 \Mem_reg[44][10]  ( .D(n3704), .CLK(clk), .Q(\Mem[44][10] ) );
  DFFPOSX1 \Mem_reg[44][9]  ( .D(n3703), .CLK(clk), .Q(\Mem[44][9] ) );
  DFFPOSX1 \Mem_reg[44][8]  ( .D(n3702), .CLK(clk), .Q(\Mem[44][8] ) );
  DFFPOSX1 \Mem_reg[44][7]  ( .D(n3701), .CLK(clk), .Q(\Mem[44][7] ) );
  DFFPOSX1 \Mem_reg[44][6]  ( .D(n3700), .CLK(clk), .Q(\Mem[44][6] ) );
  DFFPOSX1 \Mem_reg[44][5]  ( .D(n3699), .CLK(clk), .Q(\Mem[44][5] ) );
  DFFPOSX1 \Mem_reg[44][4]  ( .D(n3698), .CLK(clk), .Q(\Mem[44][4] ) );
  DFFPOSX1 \Mem_reg[44][3]  ( .D(n3697), .CLK(clk), .Q(\Mem[44][3] ) );
  DFFPOSX1 \Mem_reg[44][2]  ( .D(n3696), .CLK(clk), .Q(\Mem[44][2] ) );
  DFFPOSX1 \Mem_reg[44][1]  ( .D(n3695), .CLK(clk), .Q(\Mem[44][1] ) );
  DFFPOSX1 \Mem_reg[44][0]  ( .D(n3694), .CLK(clk), .Q(\Mem[44][0] ) );
  DFFPOSX1 \Mem_reg[43][31]  ( .D(n3693), .CLK(clk), .Q(\Mem[43][31] ) );
  DFFPOSX1 \Mem_reg[43][30]  ( .D(n3692), .CLK(clk), .Q(\Mem[43][30] ) );
  DFFPOSX1 \Mem_reg[43][29]  ( .D(n3691), .CLK(clk), .Q(\Mem[43][29] ) );
  DFFPOSX1 \Mem_reg[43][28]  ( .D(n3690), .CLK(clk), .Q(\Mem[43][28] ) );
  DFFPOSX1 \Mem_reg[43][27]  ( .D(n3689), .CLK(clk), .Q(\Mem[43][27] ) );
  DFFPOSX1 \Mem_reg[43][26]  ( .D(n3688), .CLK(clk), .Q(\Mem[43][26] ) );
  DFFPOSX1 \Mem_reg[43][25]  ( .D(n3687), .CLK(clk), .Q(\Mem[43][25] ) );
  DFFPOSX1 \Mem_reg[43][24]  ( .D(n3686), .CLK(clk), .Q(\Mem[43][24] ) );
  DFFPOSX1 \Mem_reg[43][23]  ( .D(n3685), .CLK(clk), .Q(\Mem[43][23] ) );
  DFFPOSX1 \Mem_reg[43][22]  ( .D(n3684), .CLK(clk), .Q(\Mem[43][22] ) );
  DFFPOSX1 \Mem_reg[43][21]  ( .D(n3683), .CLK(clk), .Q(\Mem[43][21] ) );
  DFFPOSX1 \Mem_reg[43][20]  ( .D(n3682), .CLK(clk), .Q(\Mem[43][20] ) );
  DFFPOSX1 \Mem_reg[43][19]  ( .D(n3681), .CLK(clk), .Q(\Mem[43][19] ) );
  DFFPOSX1 \Mem_reg[43][18]  ( .D(n3680), .CLK(clk), .Q(\Mem[43][18] ) );
  DFFPOSX1 \Mem_reg[43][17]  ( .D(n3679), .CLK(clk), .Q(\Mem[43][17] ) );
  DFFPOSX1 \Mem_reg[43][16]  ( .D(n3678), .CLK(clk), .Q(\Mem[43][16] ) );
  DFFPOSX1 \Mem_reg[43][15]  ( .D(n3677), .CLK(clk), .Q(\Mem[43][15] ) );
  DFFPOSX1 \Mem_reg[43][14]  ( .D(n3676), .CLK(clk), .Q(\Mem[43][14] ) );
  DFFPOSX1 \Mem_reg[43][13]  ( .D(n3675), .CLK(clk), .Q(\Mem[43][13] ) );
  DFFPOSX1 \Mem_reg[43][12]  ( .D(n3674), .CLK(clk), .Q(\Mem[43][12] ) );
  DFFPOSX1 \Mem_reg[43][11]  ( .D(n3673), .CLK(clk), .Q(\Mem[43][11] ) );
  DFFPOSX1 \Mem_reg[43][10]  ( .D(n3672), .CLK(clk), .Q(\Mem[43][10] ) );
  DFFPOSX1 \Mem_reg[43][9]  ( .D(n3671), .CLK(clk), .Q(\Mem[43][9] ) );
  DFFPOSX1 \Mem_reg[43][8]  ( .D(n3670), .CLK(clk), .Q(\Mem[43][8] ) );
  DFFPOSX1 \Mem_reg[43][7]  ( .D(n3669), .CLK(clk), .Q(\Mem[43][7] ) );
  DFFPOSX1 \Mem_reg[43][6]  ( .D(n3668), .CLK(clk), .Q(\Mem[43][6] ) );
  DFFPOSX1 \Mem_reg[43][5]  ( .D(n3667), .CLK(clk), .Q(\Mem[43][5] ) );
  DFFPOSX1 \Mem_reg[43][4]  ( .D(n3666), .CLK(clk), .Q(\Mem[43][4] ) );
  DFFPOSX1 \Mem_reg[43][3]  ( .D(n3665), .CLK(clk), .Q(\Mem[43][3] ) );
  DFFPOSX1 \Mem_reg[43][2]  ( .D(n3664), .CLK(clk), .Q(\Mem[43][2] ) );
  DFFPOSX1 \Mem_reg[43][1]  ( .D(n3663), .CLK(clk), .Q(\Mem[43][1] ) );
  DFFPOSX1 \Mem_reg[43][0]  ( .D(n3662), .CLK(clk), .Q(\Mem[43][0] ) );
  DFFPOSX1 \Mem_reg[42][31]  ( .D(n3661), .CLK(clk), .Q(\Mem[42][31] ) );
  DFFPOSX1 \Mem_reg[42][30]  ( .D(n3660), .CLK(clk), .Q(\Mem[42][30] ) );
  DFFPOSX1 \Mem_reg[42][29]  ( .D(n3659), .CLK(clk), .Q(\Mem[42][29] ) );
  DFFPOSX1 \Mem_reg[42][28]  ( .D(n3658), .CLK(clk), .Q(\Mem[42][28] ) );
  DFFPOSX1 \Mem_reg[42][27]  ( .D(n3657), .CLK(clk), .Q(\Mem[42][27] ) );
  DFFPOSX1 \Mem_reg[42][26]  ( .D(n3656), .CLK(clk), .Q(\Mem[42][26] ) );
  DFFPOSX1 \Mem_reg[42][25]  ( .D(n3655), .CLK(clk), .Q(\Mem[42][25] ) );
  DFFPOSX1 \Mem_reg[42][24]  ( .D(n3654), .CLK(clk), .Q(\Mem[42][24] ) );
  DFFPOSX1 \Mem_reg[42][23]  ( .D(n3653), .CLK(clk), .Q(\Mem[42][23] ) );
  DFFPOSX1 \Mem_reg[42][22]  ( .D(n3652), .CLK(clk), .Q(\Mem[42][22] ) );
  DFFPOSX1 \Mem_reg[42][21]  ( .D(n3651), .CLK(clk), .Q(\Mem[42][21] ) );
  DFFPOSX1 \Mem_reg[42][20]  ( .D(n3650), .CLK(clk), .Q(\Mem[42][20] ) );
  DFFPOSX1 \Mem_reg[42][19]  ( .D(n3649), .CLK(clk), .Q(\Mem[42][19] ) );
  DFFPOSX1 \Mem_reg[42][18]  ( .D(n3648), .CLK(clk), .Q(\Mem[42][18] ) );
  DFFPOSX1 \Mem_reg[42][17]  ( .D(n3647), .CLK(clk), .Q(\Mem[42][17] ) );
  DFFPOSX1 \Mem_reg[42][16]  ( .D(n3646), .CLK(clk), .Q(\Mem[42][16] ) );
  DFFPOSX1 \Mem_reg[42][15]  ( .D(n3645), .CLK(clk), .Q(\Mem[42][15] ) );
  DFFPOSX1 \Mem_reg[42][14]  ( .D(n3644), .CLK(clk), .Q(\Mem[42][14] ) );
  DFFPOSX1 \Mem_reg[42][13]  ( .D(n3643), .CLK(clk), .Q(\Mem[42][13] ) );
  DFFPOSX1 \Mem_reg[42][12]  ( .D(n3642), .CLK(clk), .Q(\Mem[42][12] ) );
  DFFPOSX1 \Mem_reg[42][11]  ( .D(n3641), .CLK(clk), .Q(\Mem[42][11] ) );
  DFFPOSX1 \Mem_reg[42][10]  ( .D(n3640), .CLK(clk), .Q(\Mem[42][10] ) );
  DFFPOSX1 \Mem_reg[42][9]  ( .D(n3639), .CLK(clk), .Q(\Mem[42][9] ) );
  DFFPOSX1 \Mem_reg[42][8]  ( .D(n3638), .CLK(clk), .Q(\Mem[42][8] ) );
  DFFPOSX1 \Mem_reg[42][7]  ( .D(n3637), .CLK(clk), .Q(\Mem[42][7] ) );
  DFFPOSX1 \Mem_reg[42][6]  ( .D(n3636), .CLK(clk), .Q(\Mem[42][6] ) );
  DFFPOSX1 \Mem_reg[42][5]  ( .D(n3635), .CLK(clk), .Q(\Mem[42][5] ) );
  DFFPOSX1 \Mem_reg[42][4]  ( .D(n3634), .CLK(clk), .Q(\Mem[42][4] ) );
  DFFPOSX1 \Mem_reg[42][3]  ( .D(n3633), .CLK(clk), .Q(\Mem[42][3] ) );
  DFFPOSX1 \Mem_reg[42][2]  ( .D(n3632), .CLK(clk), .Q(\Mem[42][2] ) );
  DFFPOSX1 \Mem_reg[42][1]  ( .D(n3631), .CLK(clk), .Q(\Mem[42][1] ) );
  DFFPOSX1 \Mem_reg[42][0]  ( .D(n3630), .CLK(clk), .Q(\Mem[42][0] ) );
  DFFPOSX1 \Mem_reg[41][31]  ( .D(n3629), .CLK(clk), .Q(\Mem[41][31] ) );
  DFFPOSX1 \Mem_reg[41][30]  ( .D(n3628), .CLK(clk), .Q(\Mem[41][30] ) );
  DFFPOSX1 \Mem_reg[41][29]  ( .D(n3627), .CLK(clk), .Q(\Mem[41][29] ) );
  DFFPOSX1 \Mem_reg[41][28]  ( .D(n3626), .CLK(clk), .Q(\Mem[41][28] ) );
  DFFPOSX1 \Mem_reg[41][27]  ( .D(n3625), .CLK(clk), .Q(\Mem[41][27] ) );
  DFFPOSX1 \Mem_reg[41][26]  ( .D(n3624), .CLK(clk), .Q(\Mem[41][26] ) );
  DFFPOSX1 \Mem_reg[41][25]  ( .D(n3623), .CLK(clk), .Q(\Mem[41][25] ) );
  DFFPOSX1 \Mem_reg[41][24]  ( .D(n3622), .CLK(clk), .Q(\Mem[41][24] ) );
  DFFPOSX1 \Mem_reg[41][23]  ( .D(n3621), .CLK(clk), .Q(\Mem[41][23] ) );
  DFFPOSX1 \Mem_reg[41][22]  ( .D(n3620), .CLK(clk), .Q(\Mem[41][22] ) );
  DFFPOSX1 \Mem_reg[41][21]  ( .D(n3619), .CLK(clk), .Q(\Mem[41][21] ) );
  DFFPOSX1 \Mem_reg[41][20]  ( .D(n3618), .CLK(clk), .Q(\Mem[41][20] ) );
  DFFPOSX1 \Mem_reg[41][19]  ( .D(n3617), .CLK(clk), .Q(\Mem[41][19] ) );
  DFFPOSX1 \Mem_reg[41][18]  ( .D(n3616), .CLK(clk), .Q(\Mem[41][18] ) );
  DFFPOSX1 \Mem_reg[41][17]  ( .D(n3615), .CLK(clk), .Q(\Mem[41][17] ) );
  DFFPOSX1 \Mem_reg[41][16]  ( .D(n3614), .CLK(clk), .Q(\Mem[41][16] ) );
  DFFPOSX1 \Mem_reg[41][15]  ( .D(n3613), .CLK(clk), .Q(\Mem[41][15] ) );
  DFFPOSX1 \Mem_reg[41][14]  ( .D(n3612), .CLK(clk), .Q(\Mem[41][14] ) );
  DFFPOSX1 \Mem_reg[41][13]  ( .D(n3611), .CLK(clk), .Q(\Mem[41][13] ) );
  DFFPOSX1 \Mem_reg[41][12]  ( .D(n3610), .CLK(clk), .Q(\Mem[41][12] ) );
  DFFPOSX1 \Mem_reg[41][11]  ( .D(n3609), .CLK(clk), .Q(\Mem[41][11] ) );
  DFFPOSX1 \Mem_reg[41][10]  ( .D(n3608), .CLK(clk), .Q(\Mem[41][10] ) );
  DFFPOSX1 \Mem_reg[41][9]  ( .D(n3607), .CLK(clk), .Q(\Mem[41][9] ) );
  DFFPOSX1 \Mem_reg[41][8]  ( .D(n3606), .CLK(clk), .Q(\Mem[41][8] ) );
  DFFPOSX1 \Mem_reg[41][7]  ( .D(n3605), .CLK(clk), .Q(\Mem[41][7] ) );
  DFFPOSX1 \Mem_reg[41][6]  ( .D(n3604), .CLK(clk), .Q(\Mem[41][6] ) );
  DFFPOSX1 \Mem_reg[41][5]  ( .D(n3603), .CLK(clk), .Q(\Mem[41][5] ) );
  DFFPOSX1 \Mem_reg[41][4]  ( .D(n3602), .CLK(clk), .Q(\Mem[41][4] ) );
  DFFPOSX1 \Mem_reg[41][3]  ( .D(n3601), .CLK(clk), .Q(\Mem[41][3] ) );
  DFFPOSX1 \Mem_reg[41][2]  ( .D(n3600), .CLK(clk), .Q(\Mem[41][2] ) );
  DFFPOSX1 \Mem_reg[41][1]  ( .D(n3599), .CLK(clk), .Q(\Mem[41][1] ) );
  DFFPOSX1 \Mem_reg[41][0]  ( .D(n3598), .CLK(clk), .Q(\Mem[41][0] ) );
  DFFPOSX1 \Mem_reg[40][31]  ( .D(n3597), .CLK(clk), .Q(\Mem[40][31] ) );
  DFFPOSX1 \Mem_reg[40][30]  ( .D(n3596), .CLK(clk), .Q(\Mem[40][30] ) );
  DFFPOSX1 \Mem_reg[40][29]  ( .D(n3595), .CLK(clk), .Q(\Mem[40][29] ) );
  DFFPOSX1 \Mem_reg[40][28]  ( .D(n3594), .CLK(clk), .Q(\Mem[40][28] ) );
  DFFPOSX1 \Mem_reg[40][27]  ( .D(n3593), .CLK(clk), .Q(\Mem[40][27] ) );
  DFFPOSX1 \Mem_reg[40][26]  ( .D(n3592), .CLK(clk), .Q(\Mem[40][26] ) );
  DFFPOSX1 \Mem_reg[40][25]  ( .D(n3591), .CLK(clk), .Q(\Mem[40][25] ) );
  DFFPOSX1 \Mem_reg[40][24]  ( .D(n3590), .CLK(clk), .Q(\Mem[40][24] ) );
  DFFPOSX1 \Mem_reg[40][23]  ( .D(n3589), .CLK(clk), .Q(\Mem[40][23] ) );
  DFFPOSX1 \Mem_reg[40][22]  ( .D(n3588), .CLK(clk), .Q(\Mem[40][22] ) );
  DFFPOSX1 \Mem_reg[40][21]  ( .D(n3587), .CLK(clk), .Q(\Mem[40][21] ) );
  DFFPOSX1 \Mem_reg[40][20]  ( .D(n3586), .CLK(clk), .Q(\Mem[40][20] ) );
  DFFPOSX1 \Mem_reg[40][19]  ( .D(n3585), .CLK(clk), .Q(\Mem[40][19] ) );
  DFFPOSX1 \Mem_reg[40][18]  ( .D(n3584), .CLK(clk), .Q(\Mem[40][18] ) );
  DFFPOSX1 \Mem_reg[40][17]  ( .D(n3583), .CLK(clk), .Q(\Mem[40][17] ) );
  DFFPOSX1 \Mem_reg[40][16]  ( .D(n3582), .CLK(clk), .Q(\Mem[40][16] ) );
  DFFPOSX1 \Mem_reg[40][15]  ( .D(n3581), .CLK(clk), .Q(\Mem[40][15] ) );
  DFFPOSX1 \Mem_reg[40][14]  ( .D(n3580), .CLK(clk), .Q(\Mem[40][14] ) );
  DFFPOSX1 \Mem_reg[40][13]  ( .D(n3579), .CLK(clk), .Q(\Mem[40][13] ) );
  DFFPOSX1 \Mem_reg[40][12]  ( .D(n3578), .CLK(clk), .Q(\Mem[40][12] ) );
  DFFPOSX1 \Mem_reg[40][11]  ( .D(n3577), .CLK(clk), .Q(\Mem[40][11] ) );
  DFFPOSX1 \Mem_reg[40][10]  ( .D(n3576), .CLK(clk), .Q(\Mem[40][10] ) );
  DFFPOSX1 \Mem_reg[40][9]  ( .D(n3575), .CLK(clk), .Q(\Mem[40][9] ) );
  DFFPOSX1 \Mem_reg[40][8]  ( .D(n3574), .CLK(clk), .Q(\Mem[40][8] ) );
  DFFPOSX1 \Mem_reg[40][7]  ( .D(n3573), .CLK(clk), .Q(\Mem[40][7] ) );
  DFFPOSX1 \Mem_reg[40][6]  ( .D(n3572), .CLK(clk), .Q(\Mem[40][6] ) );
  DFFPOSX1 \Mem_reg[40][5]  ( .D(n3571), .CLK(clk), .Q(\Mem[40][5] ) );
  DFFPOSX1 \Mem_reg[40][4]  ( .D(n3570), .CLK(clk), .Q(\Mem[40][4] ) );
  DFFPOSX1 \Mem_reg[40][3]  ( .D(n3569), .CLK(clk), .Q(\Mem[40][3] ) );
  DFFPOSX1 \Mem_reg[40][2]  ( .D(n3568), .CLK(clk), .Q(\Mem[40][2] ) );
  DFFPOSX1 \Mem_reg[40][1]  ( .D(n3567), .CLK(clk), .Q(\Mem[40][1] ) );
  DFFPOSX1 \Mem_reg[40][0]  ( .D(n3566), .CLK(clk), .Q(\Mem[40][0] ) );
  DFFPOSX1 \Mem_reg[39][31]  ( .D(n3565), .CLK(clk), .Q(\Mem[39][31] ) );
  DFFPOSX1 \Mem_reg[39][30]  ( .D(n3564), .CLK(clk), .Q(\Mem[39][30] ) );
  DFFPOSX1 \Mem_reg[39][29]  ( .D(n3563), .CLK(clk), .Q(\Mem[39][29] ) );
  DFFPOSX1 \Mem_reg[39][28]  ( .D(n3562), .CLK(clk), .Q(\Mem[39][28] ) );
  DFFPOSX1 \Mem_reg[39][27]  ( .D(n3561), .CLK(clk), .Q(\Mem[39][27] ) );
  DFFPOSX1 \Mem_reg[39][26]  ( .D(n3560), .CLK(clk), .Q(\Mem[39][26] ) );
  DFFPOSX1 \Mem_reg[39][25]  ( .D(n3559), .CLK(clk), .Q(\Mem[39][25] ) );
  DFFPOSX1 \Mem_reg[39][24]  ( .D(n3558), .CLK(clk), .Q(\Mem[39][24] ) );
  DFFPOSX1 \Mem_reg[39][23]  ( .D(n3557), .CLK(clk), .Q(\Mem[39][23] ) );
  DFFPOSX1 \Mem_reg[39][22]  ( .D(n3556), .CLK(clk), .Q(\Mem[39][22] ) );
  DFFPOSX1 \Mem_reg[39][21]  ( .D(n3555), .CLK(clk), .Q(\Mem[39][21] ) );
  DFFPOSX1 \Mem_reg[39][20]  ( .D(n3554), .CLK(clk), .Q(\Mem[39][20] ) );
  DFFPOSX1 \Mem_reg[39][19]  ( .D(n3553), .CLK(clk), .Q(\Mem[39][19] ) );
  DFFPOSX1 \Mem_reg[39][18]  ( .D(n3552), .CLK(clk), .Q(\Mem[39][18] ) );
  DFFPOSX1 \Mem_reg[39][17]  ( .D(n3551), .CLK(clk), .Q(\Mem[39][17] ) );
  DFFPOSX1 \Mem_reg[39][16]  ( .D(n3550), .CLK(clk), .Q(\Mem[39][16] ) );
  DFFPOSX1 \Mem_reg[39][15]  ( .D(n3549), .CLK(clk), .Q(\Mem[39][15] ) );
  DFFPOSX1 \Mem_reg[39][14]  ( .D(n3548), .CLK(clk), .Q(\Mem[39][14] ) );
  DFFPOSX1 \Mem_reg[39][13]  ( .D(n3547), .CLK(clk), .Q(\Mem[39][13] ) );
  DFFPOSX1 \Mem_reg[39][12]  ( .D(n3546), .CLK(clk), .Q(\Mem[39][12] ) );
  DFFPOSX1 \Mem_reg[39][11]  ( .D(n3545), .CLK(clk), .Q(\Mem[39][11] ) );
  DFFPOSX1 \Mem_reg[39][10]  ( .D(n3544), .CLK(clk), .Q(\Mem[39][10] ) );
  DFFPOSX1 \Mem_reg[39][9]  ( .D(n3543), .CLK(clk), .Q(\Mem[39][9] ) );
  DFFPOSX1 \Mem_reg[39][8]  ( .D(n3542), .CLK(clk), .Q(\Mem[39][8] ) );
  DFFPOSX1 \Mem_reg[39][7]  ( .D(n3541), .CLK(clk), .Q(\Mem[39][7] ) );
  DFFPOSX1 \Mem_reg[39][6]  ( .D(n3540), .CLK(clk), .Q(\Mem[39][6] ) );
  DFFPOSX1 \Mem_reg[39][5]  ( .D(n3539), .CLK(clk), .Q(\Mem[39][5] ) );
  DFFPOSX1 \Mem_reg[39][4]  ( .D(n3538), .CLK(clk), .Q(\Mem[39][4] ) );
  DFFPOSX1 \Mem_reg[39][3]  ( .D(n3537), .CLK(clk), .Q(\Mem[39][3] ) );
  DFFPOSX1 \Mem_reg[39][2]  ( .D(n3536), .CLK(clk), .Q(\Mem[39][2] ) );
  DFFPOSX1 \Mem_reg[39][1]  ( .D(n3535), .CLK(clk), .Q(\Mem[39][1] ) );
  DFFPOSX1 \Mem_reg[39][0]  ( .D(n3534), .CLK(clk), .Q(\Mem[39][0] ) );
  DFFPOSX1 \Mem_reg[38][31]  ( .D(n3533), .CLK(clk), .Q(\Mem[38][31] ) );
  DFFPOSX1 \Mem_reg[38][30]  ( .D(n3532), .CLK(clk), .Q(\Mem[38][30] ) );
  DFFPOSX1 \Mem_reg[38][29]  ( .D(n3531), .CLK(clk), .Q(\Mem[38][29] ) );
  DFFPOSX1 \Mem_reg[38][28]  ( .D(n3530), .CLK(clk), .Q(\Mem[38][28] ) );
  DFFPOSX1 \Mem_reg[38][27]  ( .D(n3529), .CLK(clk), .Q(\Mem[38][27] ) );
  DFFPOSX1 \Mem_reg[38][26]  ( .D(n3528), .CLK(clk), .Q(\Mem[38][26] ) );
  DFFPOSX1 \Mem_reg[38][25]  ( .D(n3527), .CLK(clk), .Q(\Mem[38][25] ) );
  DFFPOSX1 \Mem_reg[38][24]  ( .D(n3526), .CLK(clk), .Q(\Mem[38][24] ) );
  DFFPOSX1 \Mem_reg[38][23]  ( .D(n3525), .CLK(clk), .Q(\Mem[38][23] ) );
  DFFPOSX1 \Mem_reg[38][22]  ( .D(n3524), .CLK(clk), .Q(\Mem[38][22] ) );
  DFFPOSX1 \Mem_reg[38][21]  ( .D(n3523), .CLK(clk), .Q(\Mem[38][21] ) );
  DFFPOSX1 \Mem_reg[38][20]  ( .D(n3522), .CLK(clk), .Q(\Mem[38][20] ) );
  DFFPOSX1 \Mem_reg[38][19]  ( .D(n3521), .CLK(clk), .Q(\Mem[38][19] ) );
  DFFPOSX1 \Mem_reg[38][18]  ( .D(n3520), .CLK(clk), .Q(\Mem[38][18] ) );
  DFFPOSX1 \Mem_reg[38][17]  ( .D(n3519), .CLK(clk), .Q(\Mem[38][17] ) );
  DFFPOSX1 \Mem_reg[38][16]  ( .D(n3518), .CLK(clk), .Q(\Mem[38][16] ) );
  DFFPOSX1 \Mem_reg[38][15]  ( .D(n3517), .CLK(clk), .Q(\Mem[38][15] ) );
  DFFPOSX1 \Mem_reg[38][14]  ( .D(n3516), .CLK(clk), .Q(\Mem[38][14] ) );
  DFFPOSX1 \Mem_reg[38][13]  ( .D(n3515), .CLK(clk), .Q(\Mem[38][13] ) );
  DFFPOSX1 \Mem_reg[38][12]  ( .D(n3514), .CLK(clk), .Q(\Mem[38][12] ) );
  DFFPOSX1 \Mem_reg[38][11]  ( .D(n3513), .CLK(clk), .Q(\Mem[38][11] ) );
  DFFPOSX1 \Mem_reg[38][10]  ( .D(n3512), .CLK(clk), .Q(\Mem[38][10] ) );
  DFFPOSX1 \Mem_reg[38][9]  ( .D(n3511), .CLK(clk), .Q(\Mem[38][9] ) );
  DFFPOSX1 \Mem_reg[38][8]  ( .D(n3510), .CLK(clk), .Q(\Mem[38][8] ) );
  DFFPOSX1 \Mem_reg[38][7]  ( .D(n3509), .CLK(clk), .Q(\Mem[38][7] ) );
  DFFPOSX1 \Mem_reg[38][6]  ( .D(n3508), .CLK(clk), .Q(\Mem[38][6] ) );
  DFFPOSX1 \Mem_reg[38][5]  ( .D(n3507), .CLK(clk), .Q(\Mem[38][5] ) );
  DFFPOSX1 \Mem_reg[38][4]  ( .D(n3506), .CLK(clk), .Q(\Mem[38][4] ) );
  DFFPOSX1 \Mem_reg[38][3]  ( .D(n3505), .CLK(clk), .Q(\Mem[38][3] ) );
  DFFPOSX1 \Mem_reg[38][2]  ( .D(n3504), .CLK(clk), .Q(\Mem[38][2] ) );
  DFFPOSX1 \Mem_reg[38][1]  ( .D(n3503), .CLK(clk), .Q(\Mem[38][1] ) );
  DFFPOSX1 \Mem_reg[38][0]  ( .D(n3502), .CLK(clk), .Q(\Mem[38][0] ) );
  DFFPOSX1 \Mem_reg[37][31]  ( .D(n3501), .CLK(clk), .Q(\Mem[37][31] ) );
  DFFPOSX1 \Mem_reg[37][30]  ( .D(n3500), .CLK(clk), .Q(\Mem[37][30] ) );
  DFFPOSX1 \Mem_reg[37][29]  ( .D(n3499), .CLK(clk), .Q(\Mem[37][29] ) );
  DFFPOSX1 \Mem_reg[37][28]  ( .D(n3498), .CLK(clk), .Q(\Mem[37][28] ) );
  DFFPOSX1 \Mem_reg[37][27]  ( .D(n3497), .CLK(clk), .Q(\Mem[37][27] ) );
  DFFPOSX1 \Mem_reg[37][26]  ( .D(n3496), .CLK(clk), .Q(\Mem[37][26] ) );
  DFFPOSX1 \Mem_reg[37][25]  ( .D(n3495), .CLK(clk), .Q(\Mem[37][25] ) );
  DFFPOSX1 \Mem_reg[37][24]  ( .D(n3494), .CLK(clk), .Q(\Mem[37][24] ) );
  DFFPOSX1 \Mem_reg[37][23]  ( .D(n3493), .CLK(clk), .Q(\Mem[37][23] ) );
  DFFPOSX1 \Mem_reg[37][22]  ( .D(n3492), .CLK(clk), .Q(\Mem[37][22] ) );
  DFFPOSX1 \Mem_reg[37][21]  ( .D(n3491), .CLK(clk), .Q(\Mem[37][21] ) );
  DFFPOSX1 \Mem_reg[37][20]  ( .D(n3490), .CLK(clk), .Q(\Mem[37][20] ) );
  DFFPOSX1 \Mem_reg[37][19]  ( .D(n3489), .CLK(clk), .Q(\Mem[37][19] ) );
  DFFPOSX1 \Mem_reg[37][18]  ( .D(n3488), .CLK(clk), .Q(\Mem[37][18] ) );
  DFFPOSX1 \Mem_reg[37][17]  ( .D(n3487), .CLK(clk), .Q(\Mem[37][17] ) );
  DFFPOSX1 \Mem_reg[37][16]  ( .D(n3486), .CLK(clk), .Q(\Mem[37][16] ) );
  DFFPOSX1 \Mem_reg[37][15]  ( .D(n3485), .CLK(clk), .Q(\Mem[37][15] ) );
  DFFPOSX1 \Mem_reg[37][14]  ( .D(n3484), .CLK(clk), .Q(\Mem[37][14] ) );
  DFFPOSX1 \Mem_reg[37][13]  ( .D(n3483), .CLK(clk), .Q(\Mem[37][13] ) );
  DFFPOSX1 \Mem_reg[37][12]  ( .D(n3482), .CLK(clk), .Q(\Mem[37][12] ) );
  DFFPOSX1 \Mem_reg[37][11]  ( .D(n3481), .CLK(clk), .Q(\Mem[37][11] ) );
  DFFPOSX1 \Mem_reg[37][10]  ( .D(n3480), .CLK(clk), .Q(\Mem[37][10] ) );
  DFFPOSX1 \Mem_reg[37][9]  ( .D(n3479), .CLK(clk), .Q(\Mem[37][9] ) );
  DFFPOSX1 \Mem_reg[37][8]  ( .D(n3478), .CLK(clk), .Q(\Mem[37][8] ) );
  DFFPOSX1 \Mem_reg[37][7]  ( .D(n3477), .CLK(clk), .Q(\Mem[37][7] ) );
  DFFPOSX1 \Mem_reg[37][6]  ( .D(n3476), .CLK(clk), .Q(\Mem[37][6] ) );
  DFFPOSX1 \Mem_reg[37][5]  ( .D(n3475), .CLK(clk), .Q(\Mem[37][5] ) );
  DFFPOSX1 \Mem_reg[37][4]  ( .D(n3474), .CLK(clk), .Q(\Mem[37][4] ) );
  DFFPOSX1 \Mem_reg[37][3]  ( .D(n3473), .CLK(clk), .Q(\Mem[37][3] ) );
  DFFPOSX1 \Mem_reg[37][2]  ( .D(n3472), .CLK(clk), .Q(\Mem[37][2] ) );
  DFFPOSX1 \Mem_reg[37][1]  ( .D(n3471), .CLK(clk), .Q(\Mem[37][1] ) );
  DFFPOSX1 \Mem_reg[37][0]  ( .D(n3470), .CLK(clk), .Q(\Mem[37][0] ) );
  DFFPOSX1 \Mem_reg[36][31]  ( .D(n3469), .CLK(clk), .Q(\Mem[36][31] ) );
  DFFPOSX1 \Mem_reg[36][30]  ( .D(n3468), .CLK(clk), .Q(\Mem[36][30] ) );
  DFFPOSX1 \Mem_reg[36][29]  ( .D(n3467), .CLK(clk), .Q(\Mem[36][29] ) );
  DFFPOSX1 \Mem_reg[36][28]  ( .D(n3466), .CLK(clk), .Q(\Mem[36][28] ) );
  DFFPOSX1 \Mem_reg[36][27]  ( .D(n3465), .CLK(clk), .Q(\Mem[36][27] ) );
  DFFPOSX1 \Mem_reg[36][26]  ( .D(n3464), .CLK(clk), .Q(\Mem[36][26] ) );
  DFFPOSX1 \Mem_reg[36][25]  ( .D(n3463), .CLK(clk), .Q(\Mem[36][25] ) );
  DFFPOSX1 \Mem_reg[36][24]  ( .D(n3462), .CLK(clk), .Q(\Mem[36][24] ) );
  DFFPOSX1 \Mem_reg[36][23]  ( .D(n3461), .CLK(clk), .Q(\Mem[36][23] ) );
  DFFPOSX1 \Mem_reg[36][22]  ( .D(n3460), .CLK(clk), .Q(\Mem[36][22] ) );
  DFFPOSX1 \Mem_reg[36][21]  ( .D(n3459), .CLK(clk), .Q(\Mem[36][21] ) );
  DFFPOSX1 \Mem_reg[36][20]  ( .D(n3458), .CLK(clk), .Q(\Mem[36][20] ) );
  DFFPOSX1 \Mem_reg[36][19]  ( .D(n3457), .CLK(clk), .Q(\Mem[36][19] ) );
  DFFPOSX1 \Mem_reg[36][18]  ( .D(n3456), .CLK(clk), .Q(\Mem[36][18] ) );
  DFFPOSX1 \Mem_reg[36][17]  ( .D(n3455), .CLK(clk), .Q(\Mem[36][17] ) );
  DFFPOSX1 \Mem_reg[36][16]  ( .D(n3454), .CLK(clk), .Q(\Mem[36][16] ) );
  DFFPOSX1 \Mem_reg[36][15]  ( .D(n3453), .CLK(clk), .Q(\Mem[36][15] ) );
  DFFPOSX1 \Mem_reg[36][14]  ( .D(n3452), .CLK(clk), .Q(\Mem[36][14] ) );
  DFFPOSX1 \Mem_reg[36][13]  ( .D(n3451), .CLK(clk), .Q(\Mem[36][13] ) );
  DFFPOSX1 \Mem_reg[36][12]  ( .D(n3450), .CLK(clk), .Q(\Mem[36][12] ) );
  DFFPOSX1 \Mem_reg[36][11]  ( .D(n3449), .CLK(clk), .Q(\Mem[36][11] ) );
  DFFPOSX1 \Mem_reg[36][10]  ( .D(n3448), .CLK(clk), .Q(\Mem[36][10] ) );
  DFFPOSX1 \Mem_reg[36][9]  ( .D(n3447), .CLK(clk), .Q(\Mem[36][9] ) );
  DFFPOSX1 \Mem_reg[36][8]  ( .D(n3446), .CLK(clk), .Q(\Mem[36][8] ) );
  DFFPOSX1 \Mem_reg[36][7]  ( .D(n3445), .CLK(clk), .Q(\Mem[36][7] ) );
  DFFPOSX1 \Mem_reg[36][6]  ( .D(n3444), .CLK(clk), .Q(\Mem[36][6] ) );
  DFFPOSX1 \Mem_reg[36][5]  ( .D(n3443), .CLK(clk), .Q(\Mem[36][5] ) );
  DFFPOSX1 \Mem_reg[36][4]  ( .D(n3442), .CLK(clk), .Q(\Mem[36][4] ) );
  DFFPOSX1 \Mem_reg[36][3]  ( .D(n3441), .CLK(clk), .Q(\Mem[36][3] ) );
  DFFPOSX1 \Mem_reg[36][2]  ( .D(n3440), .CLK(clk), .Q(\Mem[36][2] ) );
  DFFPOSX1 \Mem_reg[36][1]  ( .D(n3439), .CLK(clk), .Q(\Mem[36][1] ) );
  DFFPOSX1 \Mem_reg[36][0]  ( .D(n3438), .CLK(clk), .Q(\Mem[36][0] ) );
  DFFPOSX1 \Mem_reg[35][31]  ( .D(n3437), .CLK(clk), .Q(\Mem[35][31] ) );
  DFFPOSX1 \Mem_reg[35][30]  ( .D(n3436), .CLK(clk), .Q(\Mem[35][30] ) );
  DFFPOSX1 \Mem_reg[35][29]  ( .D(n3435), .CLK(clk), .Q(\Mem[35][29] ) );
  DFFPOSX1 \Mem_reg[35][28]  ( .D(n3434), .CLK(clk), .Q(\Mem[35][28] ) );
  DFFPOSX1 \Mem_reg[35][27]  ( .D(n3433), .CLK(clk), .Q(\Mem[35][27] ) );
  DFFPOSX1 \Mem_reg[35][26]  ( .D(n3432), .CLK(clk), .Q(\Mem[35][26] ) );
  DFFPOSX1 \Mem_reg[35][25]  ( .D(n3431), .CLK(clk), .Q(\Mem[35][25] ) );
  DFFPOSX1 \Mem_reg[35][24]  ( .D(n3430), .CLK(clk), .Q(\Mem[35][24] ) );
  DFFPOSX1 \Mem_reg[35][23]  ( .D(n3429), .CLK(clk), .Q(\Mem[35][23] ) );
  DFFPOSX1 \Mem_reg[35][22]  ( .D(n3428), .CLK(clk), .Q(\Mem[35][22] ) );
  DFFPOSX1 \Mem_reg[35][21]  ( .D(n3427), .CLK(clk), .Q(\Mem[35][21] ) );
  DFFPOSX1 \Mem_reg[35][20]  ( .D(n3426), .CLK(clk), .Q(\Mem[35][20] ) );
  DFFPOSX1 \Mem_reg[35][19]  ( .D(n3425), .CLK(clk), .Q(\Mem[35][19] ) );
  DFFPOSX1 \Mem_reg[35][18]  ( .D(n3424), .CLK(clk), .Q(\Mem[35][18] ) );
  DFFPOSX1 \Mem_reg[35][17]  ( .D(n3423), .CLK(clk), .Q(\Mem[35][17] ) );
  DFFPOSX1 \Mem_reg[35][16]  ( .D(n3422), .CLK(clk), .Q(\Mem[35][16] ) );
  DFFPOSX1 \Mem_reg[35][15]  ( .D(n3421), .CLK(clk), .Q(\Mem[35][15] ) );
  DFFPOSX1 \Mem_reg[35][14]  ( .D(n3420), .CLK(clk), .Q(\Mem[35][14] ) );
  DFFPOSX1 \Mem_reg[35][13]  ( .D(n3419), .CLK(clk), .Q(\Mem[35][13] ) );
  DFFPOSX1 \Mem_reg[35][12]  ( .D(n3418), .CLK(clk), .Q(\Mem[35][12] ) );
  DFFPOSX1 \Mem_reg[35][11]  ( .D(n3417), .CLK(clk), .Q(\Mem[35][11] ) );
  DFFPOSX1 \Mem_reg[35][10]  ( .D(n3416), .CLK(clk), .Q(\Mem[35][10] ) );
  DFFPOSX1 \Mem_reg[35][9]  ( .D(n3415), .CLK(clk), .Q(\Mem[35][9] ) );
  DFFPOSX1 \Mem_reg[35][8]  ( .D(n3414), .CLK(clk), .Q(\Mem[35][8] ) );
  DFFPOSX1 \Mem_reg[35][7]  ( .D(n3413), .CLK(clk), .Q(\Mem[35][7] ) );
  DFFPOSX1 \Mem_reg[35][6]  ( .D(n3412), .CLK(clk), .Q(\Mem[35][6] ) );
  DFFPOSX1 \Mem_reg[35][5]  ( .D(n3411), .CLK(clk), .Q(\Mem[35][5] ) );
  DFFPOSX1 \Mem_reg[35][4]  ( .D(n3410), .CLK(clk), .Q(\Mem[35][4] ) );
  DFFPOSX1 \Mem_reg[35][3]  ( .D(n3409), .CLK(clk), .Q(\Mem[35][3] ) );
  DFFPOSX1 \Mem_reg[35][2]  ( .D(n3408), .CLK(clk), .Q(\Mem[35][2] ) );
  DFFPOSX1 \Mem_reg[35][1]  ( .D(n3407), .CLK(clk), .Q(\Mem[35][1] ) );
  DFFPOSX1 \Mem_reg[35][0]  ( .D(n3406), .CLK(clk), .Q(\Mem[35][0] ) );
  DFFPOSX1 \Mem_reg[34][31]  ( .D(n3405), .CLK(clk), .Q(\Mem[34][31] ) );
  DFFPOSX1 \Mem_reg[34][30]  ( .D(n3404), .CLK(clk), .Q(\Mem[34][30] ) );
  DFFPOSX1 \Mem_reg[34][29]  ( .D(n3403), .CLK(clk), .Q(\Mem[34][29] ) );
  DFFPOSX1 \Mem_reg[34][28]  ( .D(n3402), .CLK(clk), .Q(\Mem[34][28] ) );
  DFFPOSX1 \Mem_reg[34][27]  ( .D(n3401), .CLK(clk), .Q(\Mem[34][27] ) );
  DFFPOSX1 \Mem_reg[34][26]  ( .D(n3400), .CLK(clk), .Q(\Mem[34][26] ) );
  DFFPOSX1 \Mem_reg[34][25]  ( .D(n3399), .CLK(clk), .Q(\Mem[34][25] ) );
  DFFPOSX1 \Mem_reg[34][24]  ( .D(n3398), .CLK(clk), .Q(\Mem[34][24] ) );
  DFFPOSX1 \Mem_reg[34][23]  ( .D(n3397), .CLK(clk), .Q(\Mem[34][23] ) );
  DFFPOSX1 \Mem_reg[34][22]  ( .D(n3396), .CLK(clk), .Q(\Mem[34][22] ) );
  DFFPOSX1 \Mem_reg[34][21]  ( .D(n3395), .CLK(clk), .Q(\Mem[34][21] ) );
  DFFPOSX1 \Mem_reg[34][20]  ( .D(n3394), .CLK(clk), .Q(\Mem[34][20] ) );
  DFFPOSX1 \Mem_reg[34][19]  ( .D(n3393), .CLK(clk), .Q(\Mem[34][19] ) );
  DFFPOSX1 \Mem_reg[34][18]  ( .D(n3392), .CLK(clk), .Q(\Mem[34][18] ) );
  DFFPOSX1 \Mem_reg[34][17]  ( .D(n3391), .CLK(clk), .Q(\Mem[34][17] ) );
  DFFPOSX1 \Mem_reg[34][16]  ( .D(n3390), .CLK(clk), .Q(\Mem[34][16] ) );
  DFFPOSX1 \Mem_reg[34][15]  ( .D(n3389), .CLK(clk), .Q(\Mem[34][15] ) );
  DFFPOSX1 \Mem_reg[34][14]  ( .D(n3388), .CLK(clk), .Q(\Mem[34][14] ) );
  DFFPOSX1 \Mem_reg[34][13]  ( .D(n3387), .CLK(clk), .Q(\Mem[34][13] ) );
  DFFPOSX1 \Mem_reg[34][12]  ( .D(n3386), .CLK(clk), .Q(\Mem[34][12] ) );
  DFFPOSX1 \Mem_reg[34][11]  ( .D(n3385), .CLK(clk), .Q(\Mem[34][11] ) );
  DFFPOSX1 \Mem_reg[34][10]  ( .D(n3384), .CLK(clk), .Q(\Mem[34][10] ) );
  DFFPOSX1 \Mem_reg[34][9]  ( .D(n3383), .CLK(clk), .Q(\Mem[34][9] ) );
  DFFPOSX1 \Mem_reg[34][8]  ( .D(n3382), .CLK(clk), .Q(\Mem[34][8] ) );
  DFFPOSX1 \Mem_reg[34][7]  ( .D(n3381), .CLK(clk), .Q(\Mem[34][7] ) );
  DFFPOSX1 \Mem_reg[34][6]  ( .D(n3380), .CLK(clk), .Q(\Mem[34][6] ) );
  DFFPOSX1 \Mem_reg[34][5]  ( .D(n3379), .CLK(clk), .Q(\Mem[34][5] ) );
  DFFPOSX1 \Mem_reg[34][4]  ( .D(n3378), .CLK(clk), .Q(\Mem[34][4] ) );
  DFFPOSX1 \Mem_reg[34][3]  ( .D(n3377), .CLK(clk), .Q(\Mem[34][3] ) );
  DFFPOSX1 \Mem_reg[34][2]  ( .D(n3376), .CLK(clk), .Q(\Mem[34][2] ) );
  DFFPOSX1 \Mem_reg[34][1]  ( .D(n3375), .CLK(clk), .Q(\Mem[34][1] ) );
  DFFPOSX1 \Mem_reg[34][0]  ( .D(n3374), .CLK(clk), .Q(\Mem[34][0] ) );
  DFFPOSX1 \Mem_reg[33][31]  ( .D(n3373), .CLK(clk), .Q(\Mem[33][31] ) );
  DFFPOSX1 \Mem_reg[33][30]  ( .D(n3372), .CLK(clk), .Q(\Mem[33][30] ) );
  DFFPOSX1 \Mem_reg[33][29]  ( .D(n3371), .CLK(clk), .Q(\Mem[33][29] ) );
  DFFPOSX1 \Mem_reg[33][28]  ( .D(n3370), .CLK(clk), .Q(\Mem[33][28] ) );
  DFFPOSX1 \Mem_reg[33][27]  ( .D(n3369), .CLK(clk), .Q(\Mem[33][27] ) );
  DFFPOSX1 \Mem_reg[33][26]  ( .D(n3368), .CLK(clk), .Q(\Mem[33][26] ) );
  DFFPOSX1 \Mem_reg[33][25]  ( .D(n3367), .CLK(clk), .Q(\Mem[33][25] ) );
  DFFPOSX1 \Mem_reg[33][24]  ( .D(n3366), .CLK(clk), .Q(\Mem[33][24] ) );
  DFFPOSX1 \Mem_reg[33][23]  ( .D(n3365), .CLK(clk), .Q(\Mem[33][23] ) );
  DFFPOSX1 \Mem_reg[33][22]  ( .D(n3364), .CLK(clk), .Q(\Mem[33][22] ) );
  DFFPOSX1 \Mem_reg[33][21]  ( .D(n3363), .CLK(clk), .Q(\Mem[33][21] ) );
  DFFPOSX1 \Mem_reg[33][20]  ( .D(n3362), .CLK(clk), .Q(\Mem[33][20] ) );
  DFFPOSX1 \Mem_reg[33][19]  ( .D(n3361), .CLK(clk), .Q(\Mem[33][19] ) );
  DFFPOSX1 \Mem_reg[33][18]  ( .D(n3360), .CLK(clk), .Q(\Mem[33][18] ) );
  DFFPOSX1 \Mem_reg[33][17]  ( .D(n3359), .CLK(clk), .Q(\Mem[33][17] ) );
  DFFPOSX1 \Mem_reg[33][16]  ( .D(n3358), .CLK(clk), .Q(\Mem[33][16] ) );
  DFFPOSX1 \Mem_reg[33][15]  ( .D(n3357), .CLK(clk), .Q(\Mem[33][15] ) );
  DFFPOSX1 \Mem_reg[33][14]  ( .D(n3356), .CLK(clk), .Q(\Mem[33][14] ) );
  DFFPOSX1 \Mem_reg[33][13]  ( .D(n3355), .CLK(clk), .Q(\Mem[33][13] ) );
  DFFPOSX1 \Mem_reg[33][12]  ( .D(n3354), .CLK(clk), .Q(\Mem[33][12] ) );
  DFFPOSX1 \Mem_reg[33][11]  ( .D(n3353), .CLK(clk), .Q(\Mem[33][11] ) );
  DFFPOSX1 \Mem_reg[33][10]  ( .D(n3352), .CLK(clk), .Q(\Mem[33][10] ) );
  DFFPOSX1 \Mem_reg[33][9]  ( .D(n3351), .CLK(clk), .Q(\Mem[33][9] ) );
  DFFPOSX1 \Mem_reg[33][8]  ( .D(n3350), .CLK(clk), .Q(\Mem[33][8] ) );
  DFFPOSX1 \Mem_reg[33][7]  ( .D(n3349), .CLK(clk), .Q(\Mem[33][7] ) );
  DFFPOSX1 \Mem_reg[33][6]  ( .D(n3348), .CLK(clk), .Q(\Mem[33][6] ) );
  DFFPOSX1 \Mem_reg[33][5]  ( .D(n3347), .CLK(clk), .Q(\Mem[33][5] ) );
  DFFPOSX1 \Mem_reg[33][4]  ( .D(n3346), .CLK(clk), .Q(\Mem[33][4] ) );
  DFFPOSX1 \Mem_reg[33][3]  ( .D(n3345), .CLK(clk), .Q(\Mem[33][3] ) );
  DFFPOSX1 \Mem_reg[33][2]  ( .D(n3344), .CLK(clk), .Q(\Mem[33][2] ) );
  DFFPOSX1 \Mem_reg[33][1]  ( .D(n3343), .CLK(clk), .Q(\Mem[33][1] ) );
  DFFPOSX1 \Mem_reg[33][0]  ( .D(n3342), .CLK(clk), .Q(\Mem[33][0] ) );
  DFFPOSX1 \Mem_reg[32][31]  ( .D(n3341), .CLK(clk), .Q(\Mem[32][31] ) );
  DFFPOSX1 \Mem_reg[32][30]  ( .D(n3340), .CLK(clk), .Q(\Mem[32][30] ) );
  DFFPOSX1 \Mem_reg[32][29]  ( .D(n3339), .CLK(clk), .Q(\Mem[32][29] ) );
  DFFPOSX1 \Mem_reg[32][28]  ( .D(n3338), .CLK(clk), .Q(\Mem[32][28] ) );
  DFFPOSX1 \Mem_reg[32][27]  ( .D(n3337), .CLK(clk), .Q(\Mem[32][27] ) );
  DFFPOSX1 \Mem_reg[32][26]  ( .D(n3336), .CLK(clk), .Q(\Mem[32][26] ) );
  DFFPOSX1 \Mem_reg[32][25]  ( .D(n3335), .CLK(clk), .Q(\Mem[32][25] ) );
  DFFPOSX1 \Mem_reg[32][24]  ( .D(n3334), .CLK(clk), .Q(\Mem[32][24] ) );
  DFFPOSX1 \Mem_reg[32][23]  ( .D(n3333), .CLK(clk), .Q(\Mem[32][23] ) );
  DFFPOSX1 \Mem_reg[32][22]  ( .D(n3332), .CLK(clk), .Q(\Mem[32][22] ) );
  DFFPOSX1 \Mem_reg[32][21]  ( .D(n3331), .CLK(clk), .Q(\Mem[32][21] ) );
  DFFPOSX1 \Mem_reg[32][20]  ( .D(n3330), .CLK(clk), .Q(\Mem[32][20] ) );
  DFFPOSX1 \Mem_reg[32][19]  ( .D(n3329), .CLK(clk), .Q(\Mem[32][19] ) );
  DFFPOSX1 \Mem_reg[32][18]  ( .D(n3328), .CLK(clk), .Q(\Mem[32][18] ) );
  DFFPOSX1 \Mem_reg[32][17]  ( .D(n3327), .CLK(clk), .Q(\Mem[32][17] ) );
  DFFPOSX1 \Mem_reg[32][16]  ( .D(n3326), .CLK(clk), .Q(\Mem[32][16] ) );
  DFFPOSX1 \Mem_reg[32][15]  ( .D(n3325), .CLK(clk), .Q(\Mem[32][15] ) );
  DFFPOSX1 \Mem_reg[32][14]  ( .D(n3324), .CLK(clk), .Q(\Mem[32][14] ) );
  DFFPOSX1 \Mem_reg[32][13]  ( .D(n3323), .CLK(clk), .Q(\Mem[32][13] ) );
  DFFPOSX1 \Mem_reg[32][12]  ( .D(n3322), .CLK(clk), .Q(\Mem[32][12] ) );
  DFFPOSX1 \Mem_reg[32][11]  ( .D(n3321), .CLK(clk), .Q(\Mem[32][11] ) );
  DFFPOSX1 \Mem_reg[32][10]  ( .D(n3320), .CLK(clk), .Q(\Mem[32][10] ) );
  DFFPOSX1 \Mem_reg[32][9]  ( .D(n3319), .CLK(clk), .Q(\Mem[32][9] ) );
  DFFPOSX1 \Mem_reg[32][8]  ( .D(n3318), .CLK(clk), .Q(\Mem[32][8] ) );
  DFFPOSX1 \Mem_reg[32][7]  ( .D(n3317), .CLK(clk), .Q(\Mem[32][7] ) );
  DFFPOSX1 \Mem_reg[32][6]  ( .D(n3316), .CLK(clk), .Q(\Mem[32][6] ) );
  DFFPOSX1 \Mem_reg[32][5]  ( .D(n3315), .CLK(clk), .Q(\Mem[32][5] ) );
  DFFPOSX1 \Mem_reg[32][4]  ( .D(n3314), .CLK(clk), .Q(\Mem[32][4] ) );
  DFFPOSX1 \Mem_reg[32][3]  ( .D(n3313), .CLK(clk), .Q(\Mem[32][3] ) );
  DFFPOSX1 \Mem_reg[32][2]  ( .D(n3312), .CLK(clk), .Q(\Mem[32][2] ) );
  DFFPOSX1 \Mem_reg[32][1]  ( .D(n3311), .CLK(clk), .Q(\Mem[32][1] ) );
  DFFPOSX1 \Mem_reg[32][0]  ( .D(n3310), .CLK(clk), .Q(\Mem[32][0] ) );
  DFFPOSX1 \Mem_reg[31][31]  ( .D(n3309), .CLK(clk), .Q(\Mem[31][31] ) );
  DFFPOSX1 \Mem_reg[31][30]  ( .D(n3308), .CLK(clk), .Q(\Mem[31][30] ) );
  DFFPOSX1 \Mem_reg[31][29]  ( .D(n3307), .CLK(clk), .Q(\Mem[31][29] ) );
  DFFPOSX1 \Mem_reg[31][28]  ( .D(n3306), .CLK(clk), .Q(\Mem[31][28] ) );
  DFFPOSX1 \Mem_reg[31][27]  ( .D(n3305), .CLK(clk), .Q(\Mem[31][27] ) );
  DFFPOSX1 \Mem_reg[31][26]  ( .D(n3304), .CLK(clk), .Q(\Mem[31][26] ) );
  DFFPOSX1 \Mem_reg[31][25]  ( .D(n3303), .CLK(clk), .Q(\Mem[31][25] ) );
  DFFPOSX1 \Mem_reg[31][24]  ( .D(n3302), .CLK(clk), .Q(\Mem[31][24] ) );
  DFFPOSX1 \Mem_reg[31][23]  ( .D(n3301), .CLK(clk), .Q(\Mem[31][23] ) );
  DFFPOSX1 \Mem_reg[31][22]  ( .D(n3300), .CLK(clk), .Q(\Mem[31][22] ) );
  DFFPOSX1 \Mem_reg[31][21]  ( .D(n3299), .CLK(clk), .Q(\Mem[31][21] ) );
  DFFPOSX1 \Mem_reg[31][20]  ( .D(n3298), .CLK(clk), .Q(\Mem[31][20] ) );
  DFFPOSX1 \Mem_reg[31][19]  ( .D(n3297), .CLK(clk), .Q(\Mem[31][19] ) );
  DFFPOSX1 \Mem_reg[31][18]  ( .D(n3296), .CLK(clk), .Q(\Mem[31][18] ) );
  DFFPOSX1 \Mem_reg[31][17]  ( .D(n3295), .CLK(clk), .Q(\Mem[31][17] ) );
  DFFPOSX1 \Mem_reg[31][16]  ( .D(n3294), .CLK(clk), .Q(\Mem[31][16] ) );
  DFFPOSX1 \Mem_reg[31][15]  ( .D(n3293), .CLK(clk), .Q(\Mem[31][15] ) );
  DFFPOSX1 \Mem_reg[31][14]  ( .D(n3292), .CLK(clk), .Q(\Mem[31][14] ) );
  DFFPOSX1 \Mem_reg[31][13]  ( .D(n3291), .CLK(clk), .Q(\Mem[31][13] ) );
  DFFPOSX1 \Mem_reg[31][12]  ( .D(n3290), .CLK(clk), .Q(\Mem[31][12] ) );
  DFFPOSX1 \Mem_reg[31][11]  ( .D(n3289), .CLK(clk), .Q(\Mem[31][11] ) );
  DFFPOSX1 \Mem_reg[31][10]  ( .D(n3288), .CLK(clk), .Q(\Mem[31][10] ) );
  DFFPOSX1 \Mem_reg[31][9]  ( .D(n3287), .CLK(clk), .Q(\Mem[31][9] ) );
  DFFPOSX1 \Mem_reg[31][8]  ( .D(n3286), .CLK(clk), .Q(\Mem[31][8] ) );
  DFFPOSX1 \Mem_reg[31][7]  ( .D(n3285), .CLK(clk), .Q(\Mem[31][7] ) );
  DFFPOSX1 \Mem_reg[31][6]  ( .D(n3284), .CLK(clk), .Q(\Mem[31][6] ) );
  DFFPOSX1 \Mem_reg[31][5]  ( .D(n3283), .CLK(clk), .Q(\Mem[31][5] ) );
  DFFPOSX1 \Mem_reg[31][4]  ( .D(n3282), .CLK(clk), .Q(\Mem[31][4] ) );
  DFFPOSX1 \Mem_reg[31][3]  ( .D(n3281), .CLK(clk), .Q(\Mem[31][3] ) );
  DFFPOSX1 \Mem_reg[31][2]  ( .D(n3280), .CLK(clk), .Q(\Mem[31][2] ) );
  DFFPOSX1 \Mem_reg[31][1]  ( .D(n3279), .CLK(clk), .Q(\Mem[31][1] ) );
  DFFPOSX1 \Mem_reg[31][0]  ( .D(n3278), .CLK(clk), .Q(\Mem[31][0] ) );
  DFFPOSX1 \Mem_reg[30][31]  ( .D(n3277), .CLK(clk), .Q(\Mem[30][31] ) );
  DFFPOSX1 \Mem_reg[30][30]  ( .D(n3276), .CLK(clk), .Q(\Mem[30][30] ) );
  DFFPOSX1 \Mem_reg[30][29]  ( .D(n3275), .CLK(clk), .Q(\Mem[30][29] ) );
  DFFPOSX1 \Mem_reg[30][28]  ( .D(n3274), .CLK(clk), .Q(\Mem[30][28] ) );
  DFFPOSX1 \Mem_reg[30][27]  ( .D(n3273), .CLK(clk), .Q(\Mem[30][27] ) );
  DFFPOSX1 \Mem_reg[30][26]  ( .D(n3272), .CLK(clk), .Q(\Mem[30][26] ) );
  DFFPOSX1 \Mem_reg[30][25]  ( .D(n3271), .CLK(clk), .Q(\Mem[30][25] ) );
  DFFPOSX1 \Mem_reg[30][24]  ( .D(n3270), .CLK(clk), .Q(\Mem[30][24] ) );
  DFFPOSX1 \Mem_reg[30][23]  ( .D(n3269), .CLK(clk), .Q(\Mem[30][23] ) );
  DFFPOSX1 \Mem_reg[30][22]  ( .D(n3268), .CLK(clk), .Q(\Mem[30][22] ) );
  DFFPOSX1 \Mem_reg[30][21]  ( .D(n3267), .CLK(clk), .Q(\Mem[30][21] ) );
  DFFPOSX1 \Mem_reg[30][20]  ( .D(n3266), .CLK(clk), .Q(\Mem[30][20] ) );
  DFFPOSX1 \Mem_reg[30][19]  ( .D(n3265), .CLK(clk), .Q(\Mem[30][19] ) );
  DFFPOSX1 \Mem_reg[30][18]  ( .D(n3264), .CLK(clk), .Q(\Mem[30][18] ) );
  DFFPOSX1 \Mem_reg[30][17]  ( .D(n3263), .CLK(clk), .Q(\Mem[30][17] ) );
  DFFPOSX1 \Mem_reg[30][16]  ( .D(n3262), .CLK(clk), .Q(\Mem[30][16] ) );
  DFFPOSX1 \Mem_reg[30][15]  ( .D(n3261), .CLK(clk), .Q(\Mem[30][15] ) );
  DFFPOSX1 \Mem_reg[30][14]  ( .D(n3260), .CLK(clk), .Q(\Mem[30][14] ) );
  DFFPOSX1 \Mem_reg[30][13]  ( .D(n3259), .CLK(clk), .Q(\Mem[30][13] ) );
  DFFPOSX1 \Mem_reg[30][12]  ( .D(n3258), .CLK(clk), .Q(\Mem[30][12] ) );
  DFFPOSX1 \Mem_reg[30][11]  ( .D(n3257), .CLK(clk), .Q(\Mem[30][11] ) );
  DFFPOSX1 \Mem_reg[30][10]  ( .D(n3256), .CLK(clk), .Q(\Mem[30][10] ) );
  DFFPOSX1 \Mem_reg[30][9]  ( .D(n3255), .CLK(clk), .Q(\Mem[30][9] ) );
  DFFPOSX1 \Mem_reg[30][8]  ( .D(n3254), .CLK(clk), .Q(\Mem[30][8] ) );
  DFFPOSX1 \Mem_reg[30][7]  ( .D(n3253), .CLK(clk), .Q(\Mem[30][7] ) );
  DFFPOSX1 \Mem_reg[30][6]  ( .D(n3252), .CLK(clk), .Q(\Mem[30][6] ) );
  DFFPOSX1 \Mem_reg[30][5]  ( .D(n3251), .CLK(clk), .Q(\Mem[30][5] ) );
  DFFPOSX1 \Mem_reg[30][4]  ( .D(n3250), .CLK(clk), .Q(\Mem[30][4] ) );
  DFFPOSX1 \Mem_reg[30][3]  ( .D(n3249), .CLK(clk), .Q(\Mem[30][3] ) );
  DFFPOSX1 \Mem_reg[30][2]  ( .D(n3248), .CLK(clk), .Q(\Mem[30][2] ) );
  DFFPOSX1 \Mem_reg[30][1]  ( .D(n3247), .CLK(clk), .Q(\Mem[30][1] ) );
  DFFPOSX1 \Mem_reg[30][0]  ( .D(n3246), .CLK(clk), .Q(\Mem[30][0] ) );
  DFFPOSX1 \Mem_reg[29][31]  ( .D(n3245), .CLK(clk), .Q(\Mem[29][31] ) );
  DFFPOSX1 \Mem_reg[29][30]  ( .D(n3244), .CLK(clk), .Q(\Mem[29][30] ) );
  DFFPOSX1 \Mem_reg[29][29]  ( .D(n3243), .CLK(clk), .Q(\Mem[29][29] ) );
  DFFPOSX1 \Mem_reg[29][28]  ( .D(n3242), .CLK(clk), .Q(\Mem[29][28] ) );
  DFFPOSX1 \Mem_reg[29][27]  ( .D(n3241), .CLK(clk), .Q(\Mem[29][27] ) );
  DFFPOSX1 \Mem_reg[29][26]  ( .D(n3240), .CLK(clk), .Q(\Mem[29][26] ) );
  DFFPOSX1 \Mem_reg[29][25]  ( .D(n3239), .CLK(clk), .Q(\Mem[29][25] ) );
  DFFPOSX1 \Mem_reg[29][24]  ( .D(n3238), .CLK(clk), .Q(\Mem[29][24] ) );
  DFFPOSX1 \Mem_reg[29][23]  ( .D(n3237), .CLK(clk), .Q(\Mem[29][23] ) );
  DFFPOSX1 \Mem_reg[29][22]  ( .D(n3236), .CLK(clk), .Q(\Mem[29][22] ) );
  DFFPOSX1 \Mem_reg[29][21]  ( .D(n3235), .CLK(clk), .Q(\Mem[29][21] ) );
  DFFPOSX1 \Mem_reg[29][20]  ( .D(n3234), .CLK(clk), .Q(\Mem[29][20] ) );
  DFFPOSX1 \Mem_reg[29][19]  ( .D(n3233), .CLK(clk), .Q(\Mem[29][19] ) );
  DFFPOSX1 \Mem_reg[29][18]  ( .D(n3232), .CLK(clk), .Q(\Mem[29][18] ) );
  DFFPOSX1 \Mem_reg[29][17]  ( .D(n3231), .CLK(clk), .Q(\Mem[29][17] ) );
  DFFPOSX1 \Mem_reg[29][16]  ( .D(n3230), .CLK(clk), .Q(\Mem[29][16] ) );
  DFFPOSX1 \Mem_reg[29][15]  ( .D(n3229), .CLK(clk), .Q(\Mem[29][15] ) );
  DFFPOSX1 \Mem_reg[29][14]  ( .D(n3228), .CLK(clk), .Q(\Mem[29][14] ) );
  DFFPOSX1 \Mem_reg[29][13]  ( .D(n3227), .CLK(clk), .Q(\Mem[29][13] ) );
  DFFPOSX1 \Mem_reg[29][12]  ( .D(n3226), .CLK(clk), .Q(\Mem[29][12] ) );
  DFFPOSX1 \Mem_reg[29][11]  ( .D(n3225), .CLK(clk), .Q(\Mem[29][11] ) );
  DFFPOSX1 \Mem_reg[29][10]  ( .D(n3224), .CLK(clk), .Q(\Mem[29][10] ) );
  DFFPOSX1 \Mem_reg[29][9]  ( .D(n3223), .CLK(clk), .Q(\Mem[29][9] ) );
  DFFPOSX1 \Mem_reg[29][8]  ( .D(n3222), .CLK(clk), .Q(\Mem[29][8] ) );
  DFFPOSX1 \Mem_reg[29][7]  ( .D(n3221), .CLK(clk), .Q(\Mem[29][7] ) );
  DFFPOSX1 \Mem_reg[29][6]  ( .D(n3220), .CLK(clk), .Q(\Mem[29][6] ) );
  DFFPOSX1 \Mem_reg[29][5]  ( .D(n3219), .CLK(clk), .Q(\Mem[29][5] ) );
  DFFPOSX1 \Mem_reg[29][4]  ( .D(n3218), .CLK(clk), .Q(\Mem[29][4] ) );
  DFFPOSX1 \Mem_reg[29][3]  ( .D(n3217), .CLK(clk), .Q(\Mem[29][3] ) );
  DFFPOSX1 \Mem_reg[29][2]  ( .D(n3216), .CLK(clk), .Q(\Mem[29][2] ) );
  DFFPOSX1 \Mem_reg[29][1]  ( .D(n3215), .CLK(clk), .Q(\Mem[29][1] ) );
  DFFPOSX1 \Mem_reg[29][0]  ( .D(n3214), .CLK(clk), .Q(\Mem[29][0] ) );
  DFFPOSX1 \Mem_reg[28][31]  ( .D(n3213), .CLK(clk), .Q(\Mem[28][31] ) );
  DFFPOSX1 \Mem_reg[28][30]  ( .D(n3212), .CLK(clk), .Q(\Mem[28][30] ) );
  DFFPOSX1 \Mem_reg[28][29]  ( .D(n3211), .CLK(clk), .Q(\Mem[28][29] ) );
  DFFPOSX1 \Mem_reg[28][28]  ( .D(n3210), .CLK(clk), .Q(\Mem[28][28] ) );
  DFFPOSX1 \Mem_reg[28][27]  ( .D(n3209), .CLK(clk), .Q(\Mem[28][27] ) );
  DFFPOSX1 \Mem_reg[28][26]  ( .D(n3208), .CLK(clk), .Q(\Mem[28][26] ) );
  DFFPOSX1 \Mem_reg[28][25]  ( .D(n3207), .CLK(clk), .Q(\Mem[28][25] ) );
  DFFPOSX1 \Mem_reg[28][24]  ( .D(n3206), .CLK(clk), .Q(\Mem[28][24] ) );
  DFFPOSX1 \Mem_reg[28][23]  ( .D(n3205), .CLK(clk), .Q(\Mem[28][23] ) );
  DFFPOSX1 \Mem_reg[28][22]  ( .D(n3204), .CLK(clk), .Q(\Mem[28][22] ) );
  DFFPOSX1 \Mem_reg[28][21]  ( .D(n3203), .CLK(clk), .Q(\Mem[28][21] ) );
  DFFPOSX1 \Mem_reg[28][20]  ( .D(n3202), .CLK(clk), .Q(\Mem[28][20] ) );
  DFFPOSX1 \Mem_reg[28][19]  ( .D(n3201), .CLK(clk), .Q(\Mem[28][19] ) );
  DFFPOSX1 \Mem_reg[28][18]  ( .D(n3200), .CLK(clk), .Q(\Mem[28][18] ) );
  DFFPOSX1 \Mem_reg[28][17]  ( .D(n3199), .CLK(clk), .Q(\Mem[28][17] ) );
  DFFPOSX1 \Mem_reg[28][16]  ( .D(n3198), .CLK(clk), .Q(\Mem[28][16] ) );
  DFFPOSX1 \Mem_reg[28][15]  ( .D(n3197), .CLK(clk), .Q(\Mem[28][15] ) );
  DFFPOSX1 \Mem_reg[28][14]  ( .D(n3196), .CLK(clk), .Q(\Mem[28][14] ) );
  DFFPOSX1 \Mem_reg[28][13]  ( .D(n3195), .CLK(clk), .Q(\Mem[28][13] ) );
  DFFPOSX1 \Mem_reg[28][12]  ( .D(n3194), .CLK(clk), .Q(\Mem[28][12] ) );
  DFFPOSX1 \Mem_reg[28][11]  ( .D(n3193), .CLK(clk), .Q(\Mem[28][11] ) );
  DFFPOSX1 \Mem_reg[28][10]  ( .D(n3192), .CLK(clk), .Q(\Mem[28][10] ) );
  DFFPOSX1 \Mem_reg[28][9]  ( .D(n3191), .CLK(clk), .Q(\Mem[28][9] ) );
  DFFPOSX1 \Mem_reg[28][8]  ( .D(n3190), .CLK(clk), .Q(\Mem[28][8] ) );
  DFFPOSX1 \Mem_reg[28][7]  ( .D(n3189), .CLK(clk), .Q(\Mem[28][7] ) );
  DFFPOSX1 \Mem_reg[28][6]  ( .D(n3188), .CLK(clk), .Q(\Mem[28][6] ) );
  DFFPOSX1 \Mem_reg[28][5]  ( .D(n3187), .CLK(clk), .Q(\Mem[28][5] ) );
  DFFPOSX1 \Mem_reg[28][4]  ( .D(n3186), .CLK(clk), .Q(\Mem[28][4] ) );
  DFFPOSX1 \Mem_reg[28][3]  ( .D(n3185), .CLK(clk), .Q(\Mem[28][3] ) );
  DFFPOSX1 \Mem_reg[28][2]  ( .D(n3184), .CLK(clk), .Q(\Mem[28][2] ) );
  DFFPOSX1 \Mem_reg[28][1]  ( .D(n3183), .CLK(clk), .Q(\Mem[28][1] ) );
  DFFPOSX1 \Mem_reg[28][0]  ( .D(n3182), .CLK(clk), .Q(\Mem[28][0] ) );
  DFFPOSX1 \Mem_reg[27][31]  ( .D(n3181), .CLK(clk), .Q(\Mem[27][31] ) );
  DFFPOSX1 \Mem_reg[27][30]  ( .D(n3180), .CLK(clk), .Q(\Mem[27][30] ) );
  DFFPOSX1 \Mem_reg[27][29]  ( .D(n3179), .CLK(clk), .Q(\Mem[27][29] ) );
  DFFPOSX1 \Mem_reg[27][28]  ( .D(n3178), .CLK(clk), .Q(\Mem[27][28] ) );
  DFFPOSX1 \Mem_reg[27][27]  ( .D(n3177), .CLK(clk), .Q(\Mem[27][27] ) );
  DFFPOSX1 \Mem_reg[27][26]  ( .D(n3176), .CLK(clk), .Q(\Mem[27][26] ) );
  DFFPOSX1 \Mem_reg[27][25]  ( .D(n3175), .CLK(clk), .Q(\Mem[27][25] ) );
  DFFPOSX1 \Mem_reg[27][24]  ( .D(n3174), .CLK(clk), .Q(\Mem[27][24] ) );
  DFFPOSX1 \Mem_reg[27][23]  ( .D(n3173), .CLK(clk), .Q(\Mem[27][23] ) );
  DFFPOSX1 \Mem_reg[27][22]  ( .D(n3172), .CLK(clk), .Q(\Mem[27][22] ) );
  DFFPOSX1 \Mem_reg[27][21]  ( .D(n3171), .CLK(clk), .Q(\Mem[27][21] ) );
  DFFPOSX1 \Mem_reg[27][20]  ( .D(n3170), .CLK(clk), .Q(\Mem[27][20] ) );
  DFFPOSX1 \Mem_reg[27][19]  ( .D(n3169), .CLK(clk), .Q(\Mem[27][19] ) );
  DFFPOSX1 \Mem_reg[27][18]  ( .D(n3168), .CLK(clk), .Q(\Mem[27][18] ) );
  DFFPOSX1 \Mem_reg[27][17]  ( .D(n3167), .CLK(clk), .Q(\Mem[27][17] ) );
  DFFPOSX1 \Mem_reg[27][16]  ( .D(n3166), .CLK(clk), .Q(\Mem[27][16] ) );
  DFFPOSX1 \Mem_reg[27][15]  ( .D(n3165), .CLK(clk), .Q(\Mem[27][15] ) );
  DFFPOSX1 \Mem_reg[27][14]  ( .D(n3164), .CLK(clk), .Q(\Mem[27][14] ) );
  DFFPOSX1 \Mem_reg[27][13]  ( .D(n3163), .CLK(clk), .Q(\Mem[27][13] ) );
  DFFPOSX1 \Mem_reg[27][12]  ( .D(n3162), .CLK(clk), .Q(\Mem[27][12] ) );
  DFFPOSX1 \Mem_reg[27][11]  ( .D(n3161), .CLK(clk), .Q(\Mem[27][11] ) );
  DFFPOSX1 \Mem_reg[27][10]  ( .D(n3160), .CLK(clk), .Q(\Mem[27][10] ) );
  DFFPOSX1 \Mem_reg[27][9]  ( .D(n3159), .CLK(clk), .Q(\Mem[27][9] ) );
  DFFPOSX1 \Mem_reg[27][8]  ( .D(n3158), .CLK(clk), .Q(\Mem[27][8] ) );
  DFFPOSX1 \Mem_reg[27][7]  ( .D(n3157), .CLK(clk), .Q(\Mem[27][7] ) );
  DFFPOSX1 \Mem_reg[27][6]  ( .D(n3156), .CLK(clk), .Q(\Mem[27][6] ) );
  DFFPOSX1 \Mem_reg[27][5]  ( .D(n3155), .CLK(clk), .Q(\Mem[27][5] ) );
  DFFPOSX1 \Mem_reg[27][4]  ( .D(n3154), .CLK(clk), .Q(\Mem[27][4] ) );
  DFFPOSX1 \Mem_reg[27][3]  ( .D(n3153), .CLK(clk), .Q(\Mem[27][3] ) );
  DFFPOSX1 \Mem_reg[27][2]  ( .D(n3152), .CLK(clk), .Q(\Mem[27][2] ) );
  DFFPOSX1 \Mem_reg[27][1]  ( .D(n3151), .CLK(clk), .Q(\Mem[27][1] ) );
  DFFPOSX1 \Mem_reg[27][0]  ( .D(n3150), .CLK(clk), .Q(\Mem[27][0] ) );
  DFFPOSX1 \Mem_reg[26][31]  ( .D(n3149), .CLK(clk), .Q(\Mem[26][31] ) );
  DFFPOSX1 \Mem_reg[26][30]  ( .D(n3148), .CLK(clk), .Q(\Mem[26][30] ) );
  DFFPOSX1 \Mem_reg[26][29]  ( .D(n3147), .CLK(clk), .Q(\Mem[26][29] ) );
  DFFPOSX1 \Mem_reg[26][28]  ( .D(n3146), .CLK(clk), .Q(\Mem[26][28] ) );
  DFFPOSX1 \Mem_reg[26][27]  ( .D(n3145), .CLK(clk), .Q(\Mem[26][27] ) );
  DFFPOSX1 \Mem_reg[26][26]  ( .D(n3144), .CLK(clk), .Q(\Mem[26][26] ) );
  DFFPOSX1 \Mem_reg[26][25]  ( .D(n3143), .CLK(clk), .Q(\Mem[26][25] ) );
  DFFPOSX1 \Mem_reg[26][24]  ( .D(n3142), .CLK(clk), .Q(\Mem[26][24] ) );
  DFFPOSX1 \Mem_reg[26][23]  ( .D(n3141), .CLK(clk), .Q(\Mem[26][23] ) );
  DFFPOSX1 \Mem_reg[26][22]  ( .D(n3140), .CLK(clk), .Q(\Mem[26][22] ) );
  DFFPOSX1 \Mem_reg[26][21]  ( .D(n3139), .CLK(clk), .Q(\Mem[26][21] ) );
  DFFPOSX1 \Mem_reg[26][20]  ( .D(n3138), .CLK(clk), .Q(\Mem[26][20] ) );
  DFFPOSX1 \Mem_reg[26][19]  ( .D(n3137), .CLK(clk), .Q(\Mem[26][19] ) );
  DFFPOSX1 \Mem_reg[26][18]  ( .D(n3136), .CLK(clk), .Q(\Mem[26][18] ) );
  DFFPOSX1 \Mem_reg[26][17]  ( .D(n3135), .CLK(clk), .Q(\Mem[26][17] ) );
  DFFPOSX1 \Mem_reg[26][16]  ( .D(n3134), .CLK(clk), .Q(\Mem[26][16] ) );
  DFFPOSX1 \Mem_reg[26][15]  ( .D(n3133), .CLK(clk), .Q(\Mem[26][15] ) );
  DFFPOSX1 \Mem_reg[26][14]  ( .D(n3132), .CLK(clk), .Q(\Mem[26][14] ) );
  DFFPOSX1 \Mem_reg[26][13]  ( .D(n3131), .CLK(clk), .Q(\Mem[26][13] ) );
  DFFPOSX1 \Mem_reg[26][12]  ( .D(n3130), .CLK(clk), .Q(\Mem[26][12] ) );
  DFFPOSX1 \Mem_reg[26][11]  ( .D(n3129), .CLK(clk), .Q(\Mem[26][11] ) );
  DFFPOSX1 \Mem_reg[26][10]  ( .D(n3128), .CLK(clk), .Q(\Mem[26][10] ) );
  DFFPOSX1 \Mem_reg[26][9]  ( .D(n3127), .CLK(clk), .Q(\Mem[26][9] ) );
  DFFPOSX1 \Mem_reg[26][8]  ( .D(n3126), .CLK(clk), .Q(\Mem[26][8] ) );
  DFFPOSX1 \Mem_reg[26][7]  ( .D(n3125), .CLK(clk), .Q(\Mem[26][7] ) );
  DFFPOSX1 \Mem_reg[26][6]  ( .D(n3124), .CLK(clk), .Q(\Mem[26][6] ) );
  DFFPOSX1 \Mem_reg[26][5]  ( .D(n3123), .CLK(clk), .Q(\Mem[26][5] ) );
  DFFPOSX1 \Mem_reg[26][4]  ( .D(n3122), .CLK(clk), .Q(\Mem[26][4] ) );
  DFFPOSX1 \Mem_reg[26][3]  ( .D(n3121), .CLK(clk), .Q(\Mem[26][3] ) );
  DFFPOSX1 \Mem_reg[26][2]  ( .D(n3120), .CLK(clk), .Q(\Mem[26][2] ) );
  DFFPOSX1 \Mem_reg[26][1]  ( .D(n3119), .CLK(clk), .Q(\Mem[26][1] ) );
  DFFPOSX1 \Mem_reg[26][0]  ( .D(n3118), .CLK(clk), .Q(\Mem[26][0] ) );
  DFFPOSX1 \Mem_reg[25][31]  ( .D(n3117), .CLK(clk), .Q(\Mem[25][31] ) );
  DFFPOSX1 \Mem_reg[25][30]  ( .D(n3116), .CLK(clk), .Q(\Mem[25][30] ) );
  DFFPOSX1 \Mem_reg[25][29]  ( .D(n3115), .CLK(clk), .Q(\Mem[25][29] ) );
  DFFPOSX1 \Mem_reg[25][28]  ( .D(n3114), .CLK(clk), .Q(\Mem[25][28] ) );
  DFFPOSX1 \Mem_reg[25][27]  ( .D(n3113), .CLK(clk), .Q(\Mem[25][27] ) );
  DFFPOSX1 \Mem_reg[25][26]  ( .D(n3112), .CLK(clk), .Q(\Mem[25][26] ) );
  DFFPOSX1 \Mem_reg[25][25]  ( .D(n3111), .CLK(clk), .Q(\Mem[25][25] ) );
  DFFPOSX1 \Mem_reg[25][24]  ( .D(n3110), .CLK(clk), .Q(\Mem[25][24] ) );
  DFFPOSX1 \Mem_reg[25][23]  ( .D(n3109), .CLK(clk), .Q(\Mem[25][23] ) );
  DFFPOSX1 \Mem_reg[25][22]  ( .D(n3108), .CLK(clk), .Q(\Mem[25][22] ) );
  DFFPOSX1 \Mem_reg[25][21]  ( .D(n3107), .CLK(clk), .Q(\Mem[25][21] ) );
  DFFPOSX1 \Mem_reg[25][20]  ( .D(n3106), .CLK(clk), .Q(\Mem[25][20] ) );
  DFFPOSX1 \Mem_reg[25][19]  ( .D(n3105), .CLK(clk), .Q(\Mem[25][19] ) );
  DFFPOSX1 \Mem_reg[25][18]  ( .D(n3104), .CLK(clk), .Q(\Mem[25][18] ) );
  DFFPOSX1 \Mem_reg[25][17]  ( .D(n3103), .CLK(clk), .Q(\Mem[25][17] ) );
  DFFPOSX1 \Mem_reg[25][16]  ( .D(n3102), .CLK(clk), .Q(\Mem[25][16] ) );
  DFFPOSX1 \Mem_reg[25][15]  ( .D(n3101), .CLK(clk), .Q(\Mem[25][15] ) );
  DFFPOSX1 \Mem_reg[25][14]  ( .D(n3100), .CLK(clk), .Q(\Mem[25][14] ) );
  DFFPOSX1 \Mem_reg[25][13]  ( .D(n3099), .CLK(clk), .Q(\Mem[25][13] ) );
  DFFPOSX1 \Mem_reg[25][12]  ( .D(n3098), .CLK(clk), .Q(\Mem[25][12] ) );
  DFFPOSX1 \Mem_reg[25][11]  ( .D(n3097), .CLK(clk), .Q(\Mem[25][11] ) );
  DFFPOSX1 \Mem_reg[25][10]  ( .D(n3096), .CLK(clk), .Q(\Mem[25][10] ) );
  DFFPOSX1 \Mem_reg[25][9]  ( .D(n3095), .CLK(clk), .Q(\Mem[25][9] ) );
  DFFPOSX1 \Mem_reg[25][8]  ( .D(n3094), .CLK(clk), .Q(\Mem[25][8] ) );
  DFFPOSX1 \Mem_reg[25][7]  ( .D(n3093), .CLK(clk), .Q(\Mem[25][7] ) );
  DFFPOSX1 \Mem_reg[25][6]  ( .D(n3092), .CLK(clk), .Q(\Mem[25][6] ) );
  DFFPOSX1 \Mem_reg[25][5]  ( .D(n3091), .CLK(clk), .Q(\Mem[25][5] ) );
  DFFPOSX1 \Mem_reg[25][4]  ( .D(n3090), .CLK(clk), .Q(\Mem[25][4] ) );
  DFFPOSX1 \Mem_reg[25][3]  ( .D(n3089), .CLK(clk), .Q(\Mem[25][3] ) );
  DFFPOSX1 \Mem_reg[25][2]  ( .D(n3088), .CLK(clk), .Q(\Mem[25][2] ) );
  DFFPOSX1 \Mem_reg[25][1]  ( .D(n3087), .CLK(clk), .Q(\Mem[25][1] ) );
  DFFPOSX1 \Mem_reg[25][0]  ( .D(n3086), .CLK(clk), .Q(\Mem[25][0] ) );
  DFFPOSX1 \Mem_reg[24][31]  ( .D(n3085), .CLK(clk), .Q(\Mem[24][31] ) );
  DFFPOSX1 \Mem_reg[24][30]  ( .D(n3084), .CLK(clk), .Q(\Mem[24][30] ) );
  DFFPOSX1 \Mem_reg[24][29]  ( .D(n3083), .CLK(clk), .Q(\Mem[24][29] ) );
  DFFPOSX1 \Mem_reg[24][28]  ( .D(n3082), .CLK(clk), .Q(\Mem[24][28] ) );
  DFFPOSX1 \Mem_reg[24][27]  ( .D(n3081), .CLK(clk), .Q(\Mem[24][27] ) );
  DFFPOSX1 \Mem_reg[24][26]  ( .D(n3080), .CLK(clk), .Q(\Mem[24][26] ) );
  DFFPOSX1 \Mem_reg[24][25]  ( .D(n3079), .CLK(clk), .Q(\Mem[24][25] ) );
  DFFPOSX1 \Mem_reg[24][24]  ( .D(n3078), .CLK(clk), .Q(\Mem[24][24] ) );
  DFFPOSX1 \Mem_reg[24][23]  ( .D(n3077), .CLK(clk), .Q(\Mem[24][23] ) );
  DFFPOSX1 \Mem_reg[24][22]  ( .D(n3076), .CLK(clk), .Q(\Mem[24][22] ) );
  DFFPOSX1 \Mem_reg[24][21]  ( .D(n3075), .CLK(clk), .Q(\Mem[24][21] ) );
  DFFPOSX1 \Mem_reg[24][20]  ( .D(n3074), .CLK(clk), .Q(\Mem[24][20] ) );
  DFFPOSX1 \Mem_reg[24][19]  ( .D(n3073), .CLK(clk), .Q(\Mem[24][19] ) );
  DFFPOSX1 \Mem_reg[24][18]  ( .D(n3072), .CLK(clk), .Q(\Mem[24][18] ) );
  DFFPOSX1 \Mem_reg[24][17]  ( .D(n3071), .CLK(clk), .Q(\Mem[24][17] ) );
  DFFPOSX1 \Mem_reg[24][16]  ( .D(n3070), .CLK(clk), .Q(\Mem[24][16] ) );
  DFFPOSX1 \Mem_reg[24][15]  ( .D(n3069), .CLK(clk), .Q(\Mem[24][15] ) );
  DFFPOSX1 \Mem_reg[24][14]  ( .D(n3068), .CLK(clk), .Q(\Mem[24][14] ) );
  DFFPOSX1 \Mem_reg[24][13]  ( .D(n3067), .CLK(clk), .Q(\Mem[24][13] ) );
  DFFPOSX1 \Mem_reg[24][12]  ( .D(n3066), .CLK(clk), .Q(\Mem[24][12] ) );
  DFFPOSX1 \Mem_reg[24][11]  ( .D(n3065), .CLK(clk), .Q(\Mem[24][11] ) );
  DFFPOSX1 \Mem_reg[24][10]  ( .D(n3064), .CLK(clk), .Q(\Mem[24][10] ) );
  DFFPOSX1 \Mem_reg[24][9]  ( .D(n3063), .CLK(clk), .Q(\Mem[24][9] ) );
  DFFPOSX1 \Mem_reg[24][8]  ( .D(n3062), .CLK(clk), .Q(\Mem[24][8] ) );
  DFFPOSX1 \Mem_reg[24][7]  ( .D(n3061), .CLK(clk), .Q(\Mem[24][7] ) );
  DFFPOSX1 \Mem_reg[24][6]  ( .D(n3060), .CLK(clk), .Q(\Mem[24][6] ) );
  DFFPOSX1 \Mem_reg[24][5]  ( .D(n3059), .CLK(clk), .Q(\Mem[24][5] ) );
  DFFPOSX1 \Mem_reg[24][4]  ( .D(n3058), .CLK(clk), .Q(\Mem[24][4] ) );
  DFFPOSX1 \Mem_reg[24][3]  ( .D(n3057), .CLK(clk), .Q(\Mem[24][3] ) );
  DFFPOSX1 \Mem_reg[24][2]  ( .D(n3056), .CLK(clk), .Q(\Mem[24][2] ) );
  DFFPOSX1 \Mem_reg[24][1]  ( .D(n3055), .CLK(clk), .Q(\Mem[24][1] ) );
  DFFPOSX1 \Mem_reg[24][0]  ( .D(n3054), .CLK(clk), .Q(\Mem[24][0] ) );
  DFFPOSX1 \Mem_reg[23][31]  ( .D(n3053), .CLK(clk), .Q(\Mem[23][31] ) );
  DFFPOSX1 \Mem_reg[23][30]  ( .D(n3052), .CLK(clk), .Q(\Mem[23][30] ) );
  DFFPOSX1 \Mem_reg[23][29]  ( .D(n3051), .CLK(clk), .Q(\Mem[23][29] ) );
  DFFPOSX1 \Mem_reg[23][28]  ( .D(n3050), .CLK(clk), .Q(\Mem[23][28] ) );
  DFFPOSX1 \Mem_reg[23][27]  ( .D(n3049), .CLK(clk), .Q(\Mem[23][27] ) );
  DFFPOSX1 \Mem_reg[23][26]  ( .D(n3048), .CLK(clk), .Q(\Mem[23][26] ) );
  DFFPOSX1 \Mem_reg[23][25]  ( .D(n3047), .CLK(clk), .Q(\Mem[23][25] ) );
  DFFPOSX1 \Mem_reg[23][24]  ( .D(n3046), .CLK(clk), .Q(\Mem[23][24] ) );
  DFFPOSX1 \Mem_reg[23][23]  ( .D(n3045), .CLK(clk), .Q(\Mem[23][23] ) );
  DFFPOSX1 \Mem_reg[23][22]  ( .D(n3044), .CLK(clk), .Q(\Mem[23][22] ) );
  DFFPOSX1 \Mem_reg[23][21]  ( .D(n3043), .CLK(clk), .Q(\Mem[23][21] ) );
  DFFPOSX1 \Mem_reg[23][20]  ( .D(n3042), .CLK(clk), .Q(\Mem[23][20] ) );
  DFFPOSX1 \Mem_reg[23][19]  ( .D(n3041), .CLK(clk), .Q(\Mem[23][19] ) );
  DFFPOSX1 \Mem_reg[23][18]  ( .D(n3040), .CLK(clk), .Q(\Mem[23][18] ) );
  DFFPOSX1 \Mem_reg[23][17]  ( .D(n3039), .CLK(clk), .Q(\Mem[23][17] ) );
  DFFPOSX1 \Mem_reg[23][16]  ( .D(n3038), .CLK(clk), .Q(\Mem[23][16] ) );
  DFFPOSX1 \Mem_reg[23][15]  ( .D(n3037), .CLK(clk), .Q(\Mem[23][15] ) );
  DFFPOSX1 \Mem_reg[23][14]  ( .D(n3036), .CLK(clk), .Q(\Mem[23][14] ) );
  DFFPOSX1 \Mem_reg[23][13]  ( .D(n3035), .CLK(clk), .Q(\Mem[23][13] ) );
  DFFPOSX1 \Mem_reg[23][12]  ( .D(n3034), .CLK(clk), .Q(\Mem[23][12] ) );
  DFFPOSX1 \Mem_reg[23][11]  ( .D(n3033), .CLK(clk), .Q(\Mem[23][11] ) );
  DFFPOSX1 \Mem_reg[23][10]  ( .D(n3032), .CLK(clk), .Q(\Mem[23][10] ) );
  DFFPOSX1 \Mem_reg[23][9]  ( .D(n3031), .CLK(clk), .Q(\Mem[23][9] ) );
  DFFPOSX1 \Mem_reg[23][8]  ( .D(n3030), .CLK(clk), .Q(\Mem[23][8] ) );
  DFFPOSX1 \Mem_reg[23][7]  ( .D(n3029), .CLK(clk), .Q(\Mem[23][7] ) );
  DFFPOSX1 \Mem_reg[23][6]  ( .D(n3028), .CLK(clk), .Q(\Mem[23][6] ) );
  DFFPOSX1 \Mem_reg[23][5]  ( .D(n3027), .CLK(clk), .Q(\Mem[23][5] ) );
  DFFPOSX1 \Mem_reg[23][4]  ( .D(n3026), .CLK(clk), .Q(\Mem[23][4] ) );
  DFFPOSX1 \Mem_reg[23][3]  ( .D(n3025), .CLK(clk), .Q(\Mem[23][3] ) );
  DFFPOSX1 \Mem_reg[23][2]  ( .D(n3024), .CLK(clk), .Q(\Mem[23][2] ) );
  DFFPOSX1 \Mem_reg[23][1]  ( .D(n3023), .CLK(clk), .Q(\Mem[23][1] ) );
  DFFPOSX1 \Mem_reg[23][0]  ( .D(n3022), .CLK(clk), .Q(\Mem[23][0] ) );
  DFFPOSX1 \Mem_reg[22][31]  ( .D(n3021), .CLK(clk), .Q(\Mem[22][31] ) );
  DFFPOSX1 \Mem_reg[22][30]  ( .D(n3020), .CLK(clk), .Q(\Mem[22][30] ) );
  DFFPOSX1 \Mem_reg[22][29]  ( .D(n3019), .CLK(clk), .Q(\Mem[22][29] ) );
  DFFPOSX1 \Mem_reg[22][28]  ( .D(n3018), .CLK(clk), .Q(\Mem[22][28] ) );
  DFFPOSX1 \Mem_reg[22][27]  ( .D(n3017), .CLK(clk), .Q(\Mem[22][27] ) );
  DFFPOSX1 \Mem_reg[22][26]  ( .D(n3016), .CLK(clk), .Q(\Mem[22][26] ) );
  DFFPOSX1 \Mem_reg[22][25]  ( .D(n3015), .CLK(clk), .Q(\Mem[22][25] ) );
  DFFPOSX1 \Mem_reg[22][24]  ( .D(n3014), .CLK(clk), .Q(\Mem[22][24] ) );
  DFFPOSX1 \Mem_reg[22][23]  ( .D(n3013), .CLK(clk), .Q(\Mem[22][23] ) );
  DFFPOSX1 \Mem_reg[22][22]  ( .D(n3012), .CLK(clk), .Q(\Mem[22][22] ) );
  DFFPOSX1 \Mem_reg[22][21]  ( .D(n3011), .CLK(clk), .Q(\Mem[22][21] ) );
  DFFPOSX1 \Mem_reg[22][20]  ( .D(n3010), .CLK(clk), .Q(\Mem[22][20] ) );
  DFFPOSX1 \Mem_reg[22][19]  ( .D(n3009), .CLK(clk), .Q(\Mem[22][19] ) );
  DFFPOSX1 \Mem_reg[22][18]  ( .D(n3008), .CLK(clk), .Q(\Mem[22][18] ) );
  DFFPOSX1 \Mem_reg[22][17]  ( .D(n3007), .CLK(clk), .Q(\Mem[22][17] ) );
  DFFPOSX1 \Mem_reg[22][16]  ( .D(n3006), .CLK(clk), .Q(\Mem[22][16] ) );
  DFFPOSX1 \Mem_reg[22][15]  ( .D(n3005), .CLK(clk), .Q(\Mem[22][15] ) );
  DFFPOSX1 \Mem_reg[22][14]  ( .D(n3004), .CLK(clk), .Q(\Mem[22][14] ) );
  DFFPOSX1 \Mem_reg[22][13]  ( .D(n3003), .CLK(clk), .Q(\Mem[22][13] ) );
  DFFPOSX1 \Mem_reg[22][12]  ( .D(n3002), .CLK(clk), .Q(\Mem[22][12] ) );
  DFFPOSX1 \Mem_reg[22][11]  ( .D(n3001), .CLK(clk), .Q(\Mem[22][11] ) );
  DFFPOSX1 \Mem_reg[22][10]  ( .D(n3000), .CLK(clk), .Q(\Mem[22][10] ) );
  DFFPOSX1 \Mem_reg[22][9]  ( .D(n2999), .CLK(clk), .Q(\Mem[22][9] ) );
  DFFPOSX1 \Mem_reg[22][8]  ( .D(n2998), .CLK(clk), .Q(\Mem[22][8] ) );
  DFFPOSX1 \Mem_reg[22][7]  ( .D(n2997), .CLK(clk), .Q(\Mem[22][7] ) );
  DFFPOSX1 \Mem_reg[22][6]  ( .D(n2996), .CLK(clk), .Q(\Mem[22][6] ) );
  DFFPOSX1 \Mem_reg[22][5]  ( .D(n2995), .CLK(clk), .Q(\Mem[22][5] ) );
  DFFPOSX1 \Mem_reg[22][4]  ( .D(n2994), .CLK(clk), .Q(\Mem[22][4] ) );
  DFFPOSX1 \Mem_reg[22][3]  ( .D(n2993), .CLK(clk), .Q(\Mem[22][3] ) );
  DFFPOSX1 \Mem_reg[22][2]  ( .D(n2992), .CLK(clk), .Q(\Mem[22][2] ) );
  DFFPOSX1 \Mem_reg[22][1]  ( .D(n2991), .CLK(clk), .Q(\Mem[22][1] ) );
  DFFPOSX1 \Mem_reg[22][0]  ( .D(n2990), .CLK(clk), .Q(\Mem[22][0] ) );
  DFFPOSX1 \Mem_reg[21][31]  ( .D(n2989), .CLK(clk), .Q(\Mem[21][31] ) );
  DFFPOSX1 \Mem_reg[21][30]  ( .D(n2988), .CLK(clk), .Q(\Mem[21][30] ) );
  DFFPOSX1 \Mem_reg[21][29]  ( .D(n2987), .CLK(clk), .Q(\Mem[21][29] ) );
  DFFPOSX1 \Mem_reg[21][28]  ( .D(n2986), .CLK(clk), .Q(\Mem[21][28] ) );
  DFFPOSX1 \Mem_reg[21][27]  ( .D(n2985), .CLK(clk), .Q(\Mem[21][27] ) );
  DFFPOSX1 \Mem_reg[21][26]  ( .D(n2984), .CLK(clk), .Q(\Mem[21][26] ) );
  DFFPOSX1 \Mem_reg[21][25]  ( .D(n2983), .CLK(clk), .Q(\Mem[21][25] ) );
  DFFPOSX1 \Mem_reg[21][24]  ( .D(n2982), .CLK(clk), .Q(\Mem[21][24] ) );
  DFFPOSX1 \Mem_reg[21][23]  ( .D(n2981), .CLK(clk), .Q(\Mem[21][23] ) );
  DFFPOSX1 \Mem_reg[21][22]  ( .D(n2980), .CLK(clk), .Q(\Mem[21][22] ) );
  DFFPOSX1 \Mem_reg[21][21]  ( .D(n2979), .CLK(clk), .Q(\Mem[21][21] ) );
  DFFPOSX1 \Mem_reg[21][20]  ( .D(n2978), .CLK(clk), .Q(\Mem[21][20] ) );
  DFFPOSX1 \Mem_reg[21][19]  ( .D(n2977), .CLK(clk), .Q(\Mem[21][19] ) );
  DFFPOSX1 \Mem_reg[21][18]  ( .D(n2976), .CLK(clk), .Q(\Mem[21][18] ) );
  DFFPOSX1 \Mem_reg[21][17]  ( .D(n2975), .CLK(clk), .Q(\Mem[21][17] ) );
  DFFPOSX1 \Mem_reg[21][16]  ( .D(n2974), .CLK(clk), .Q(\Mem[21][16] ) );
  DFFPOSX1 \Mem_reg[21][15]  ( .D(n2973), .CLK(clk), .Q(\Mem[21][15] ) );
  DFFPOSX1 \Mem_reg[21][14]  ( .D(n2972), .CLK(clk), .Q(\Mem[21][14] ) );
  DFFPOSX1 \Mem_reg[21][13]  ( .D(n2971), .CLK(clk), .Q(\Mem[21][13] ) );
  DFFPOSX1 \Mem_reg[21][12]  ( .D(n2970), .CLK(clk), .Q(\Mem[21][12] ) );
  DFFPOSX1 \Mem_reg[21][11]  ( .D(n2969), .CLK(clk), .Q(\Mem[21][11] ) );
  DFFPOSX1 \Mem_reg[21][10]  ( .D(n2968), .CLK(clk), .Q(\Mem[21][10] ) );
  DFFPOSX1 \Mem_reg[21][9]  ( .D(n2967), .CLK(clk), .Q(\Mem[21][9] ) );
  DFFPOSX1 \Mem_reg[21][8]  ( .D(n2966), .CLK(clk), .Q(\Mem[21][8] ) );
  DFFPOSX1 \Mem_reg[21][7]  ( .D(n2965), .CLK(clk), .Q(\Mem[21][7] ) );
  DFFPOSX1 \Mem_reg[21][6]  ( .D(n2964), .CLK(clk), .Q(\Mem[21][6] ) );
  DFFPOSX1 \Mem_reg[21][5]  ( .D(n2963), .CLK(clk), .Q(\Mem[21][5] ) );
  DFFPOSX1 \Mem_reg[21][4]  ( .D(n2962), .CLK(clk), .Q(\Mem[21][4] ) );
  DFFPOSX1 \Mem_reg[21][3]  ( .D(n2961), .CLK(clk), .Q(\Mem[21][3] ) );
  DFFPOSX1 \Mem_reg[21][2]  ( .D(n2960), .CLK(clk), .Q(\Mem[21][2] ) );
  DFFPOSX1 \Mem_reg[21][1]  ( .D(n2959), .CLK(clk), .Q(\Mem[21][1] ) );
  DFFPOSX1 \Mem_reg[21][0]  ( .D(n2958), .CLK(clk), .Q(\Mem[21][0] ) );
  DFFPOSX1 \Mem_reg[20][31]  ( .D(n2957), .CLK(clk), .Q(\Mem[20][31] ) );
  DFFPOSX1 \Mem_reg[20][30]  ( .D(n2956), .CLK(clk), .Q(\Mem[20][30] ) );
  DFFPOSX1 \Mem_reg[20][29]  ( .D(n2955), .CLK(clk), .Q(\Mem[20][29] ) );
  DFFPOSX1 \Mem_reg[20][28]  ( .D(n2954), .CLK(clk), .Q(\Mem[20][28] ) );
  DFFPOSX1 \Mem_reg[20][27]  ( .D(n2953), .CLK(clk), .Q(\Mem[20][27] ) );
  DFFPOSX1 \Mem_reg[20][26]  ( .D(n2952), .CLK(clk), .Q(\Mem[20][26] ) );
  DFFPOSX1 \Mem_reg[20][25]  ( .D(n2951), .CLK(clk), .Q(\Mem[20][25] ) );
  DFFPOSX1 \Mem_reg[20][24]  ( .D(n2950), .CLK(clk), .Q(\Mem[20][24] ) );
  DFFPOSX1 \Mem_reg[20][23]  ( .D(n2949), .CLK(clk), .Q(\Mem[20][23] ) );
  DFFPOSX1 \Mem_reg[20][22]  ( .D(n2948), .CLK(clk), .Q(\Mem[20][22] ) );
  DFFPOSX1 \Mem_reg[20][21]  ( .D(n2947), .CLK(clk), .Q(\Mem[20][21] ) );
  DFFPOSX1 \Mem_reg[20][20]  ( .D(n2946), .CLK(clk), .Q(\Mem[20][20] ) );
  DFFPOSX1 \Mem_reg[20][19]  ( .D(n2945), .CLK(clk), .Q(\Mem[20][19] ) );
  DFFPOSX1 \Mem_reg[20][18]  ( .D(n2944), .CLK(clk), .Q(\Mem[20][18] ) );
  DFFPOSX1 \Mem_reg[20][17]  ( .D(n2943), .CLK(clk), .Q(\Mem[20][17] ) );
  DFFPOSX1 \Mem_reg[20][16]  ( .D(n2942), .CLK(clk), .Q(\Mem[20][16] ) );
  DFFPOSX1 \Mem_reg[20][15]  ( .D(n2941), .CLK(clk), .Q(\Mem[20][15] ) );
  DFFPOSX1 \Mem_reg[20][14]  ( .D(n2940), .CLK(clk), .Q(\Mem[20][14] ) );
  DFFPOSX1 \Mem_reg[20][13]  ( .D(n2939), .CLK(clk), .Q(\Mem[20][13] ) );
  DFFPOSX1 \Mem_reg[20][12]  ( .D(n2938), .CLK(clk), .Q(\Mem[20][12] ) );
  DFFPOSX1 \Mem_reg[20][11]  ( .D(n2937), .CLK(clk), .Q(\Mem[20][11] ) );
  DFFPOSX1 \Mem_reg[20][10]  ( .D(n2936), .CLK(clk), .Q(\Mem[20][10] ) );
  DFFPOSX1 \Mem_reg[20][9]  ( .D(n2935), .CLK(clk), .Q(\Mem[20][9] ) );
  DFFPOSX1 \Mem_reg[20][8]  ( .D(n2934), .CLK(clk), .Q(\Mem[20][8] ) );
  DFFPOSX1 \Mem_reg[20][7]  ( .D(n2933), .CLK(clk), .Q(\Mem[20][7] ) );
  DFFPOSX1 \Mem_reg[20][6]  ( .D(n2932), .CLK(clk), .Q(\Mem[20][6] ) );
  DFFPOSX1 \Mem_reg[20][5]  ( .D(n2931), .CLK(clk), .Q(\Mem[20][5] ) );
  DFFPOSX1 \Mem_reg[20][4]  ( .D(n2930), .CLK(clk), .Q(\Mem[20][4] ) );
  DFFPOSX1 \Mem_reg[20][3]  ( .D(n2929), .CLK(clk), .Q(\Mem[20][3] ) );
  DFFPOSX1 \Mem_reg[20][2]  ( .D(n2928), .CLK(clk), .Q(\Mem[20][2] ) );
  DFFPOSX1 \Mem_reg[20][1]  ( .D(n2927), .CLK(clk), .Q(\Mem[20][1] ) );
  DFFPOSX1 \Mem_reg[20][0]  ( .D(n2926), .CLK(clk), .Q(\Mem[20][0] ) );
  DFFPOSX1 \Mem_reg[19][31]  ( .D(n2925), .CLK(clk), .Q(\Mem[19][31] ) );
  DFFPOSX1 \Mem_reg[19][30]  ( .D(n2924), .CLK(clk), .Q(\Mem[19][30] ) );
  DFFPOSX1 \Mem_reg[19][29]  ( .D(n2923), .CLK(clk), .Q(\Mem[19][29] ) );
  DFFPOSX1 \Mem_reg[19][28]  ( .D(n2922), .CLK(clk), .Q(\Mem[19][28] ) );
  DFFPOSX1 \Mem_reg[19][27]  ( .D(n2921), .CLK(clk), .Q(\Mem[19][27] ) );
  DFFPOSX1 \Mem_reg[19][26]  ( .D(n2920), .CLK(clk), .Q(\Mem[19][26] ) );
  DFFPOSX1 \Mem_reg[19][25]  ( .D(n2919), .CLK(clk), .Q(\Mem[19][25] ) );
  DFFPOSX1 \Mem_reg[19][24]  ( .D(n2918), .CLK(clk), .Q(\Mem[19][24] ) );
  DFFPOSX1 \Mem_reg[19][23]  ( .D(n2917), .CLK(clk), .Q(\Mem[19][23] ) );
  DFFPOSX1 \Mem_reg[19][22]  ( .D(n2916), .CLK(clk), .Q(\Mem[19][22] ) );
  DFFPOSX1 \Mem_reg[19][21]  ( .D(n2915), .CLK(clk), .Q(\Mem[19][21] ) );
  DFFPOSX1 \Mem_reg[19][20]  ( .D(n2914), .CLK(clk), .Q(\Mem[19][20] ) );
  DFFPOSX1 \Mem_reg[19][19]  ( .D(n2913), .CLK(clk), .Q(\Mem[19][19] ) );
  DFFPOSX1 \Mem_reg[19][18]  ( .D(n2912), .CLK(clk), .Q(\Mem[19][18] ) );
  DFFPOSX1 \Mem_reg[19][17]  ( .D(n2911), .CLK(clk), .Q(\Mem[19][17] ) );
  DFFPOSX1 \Mem_reg[19][16]  ( .D(n2910), .CLK(clk), .Q(\Mem[19][16] ) );
  DFFPOSX1 \Mem_reg[19][15]  ( .D(n2909), .CLK(clk), .Q(\Mem[19][15] ) );
  DFFPOSX1 \Mem_reg[19][14]  ( .D(n2908), .CLK(clk), .Q(\Mem[19][14] ) );
  DFFPOSX1 \Mem_reg[19][13]  ( .D(n2907), .CLK(clk), .Q(\Mem[19][13] ) );
  DFFPOSX1 \Mem_reg[19][12]  ( .D(n2906), .CLK(clk), .Q(\Mem[19][12] ) );
  DFFPOSX1 \Mem_reg[19][11]  ( .D(n2905), .CLK(clk), .Q(\Mem[19][11] ) );
  DFFPOSX1 \Mem_reg[19][10]  ( .D(n2904), .CLK(clk), .Q(\Mem[19][10] ) );
  DFFPOSX1 \Mem_reg[19][9]  ( .D(n2903), .CLK(clk), .Q(\Mem[19][9] ) );
  DFFPOSX1 \Mem_reg[19][8]  ( .D(n2902), .CLK(clk), .Q(\Mem[19][8] ) );
  DFFPOSX1 \Mem_reg[19][7]  ( .D(n2901), .CLK(clk), .Q(\Mem[19][7] ) );
  DFFPOSX1 \Mem_reg[19][6]  ( .D(n2900), .CLK(clk), .Q(\Mem[19][6] ) );
  DFFPOSX1 \Mem_reg[19][5]  ( .D(n2899), .CLK(clk), .Q(\Mem[19][5] ) );
  DFFPOSX1 \Mem_reg[19][4]  ( .D(n2898), .CLK(clk), .Q(\Mem[19][4] ) );
  DFFPOSX1 \Mem_reg[19][3]  ( .D(n2897), .CLK(clk), .Q(\Mem[19][3] ) );
  DFFPOSX1 \Mem_reg[19][2]  ( .D(n2896), .CLK(clk), .Q(\Mem[19][2] ) );
  DFFPOSX1 \Mem_reg[19][1]  ( .D(n2895), .CLK(clk), .Q(\Mem[19][1] ) );
  DFFPOSX1 \Mem_reg[19][0]  ( .D(n2894), .CLK(clk), .Q(\Mem[19][0] ) );
  DFFPOSX1 \Mem_reg[18][31]  ( .D(n2893), .CLK(clk), .Q(\Mem[18][31] ) );
  DFFPOSX1 \Mem_reg[18][30]  ( .D(n2892), .CLK(clk), .Q(\Mem[18][30] ) );
  DFFPOSX1 \Mem_reg[18][29]  ( .D(n2891), .CLK(clk), .Q(\Mem[18][29] ) );
  DFFPOSX1 \Mem_reg[18][28]  ( .D(n2890), .CLK(clk), .Q(\Mem[18][28] ) );
  DFFPOSX1 \Mem_reg[18][27]  ( .D(n2889), .CLK(clk), .Q(\Mem[18][27] ) );
  DFFPOSX1 \Mem_reg[18][26]  ( .D(n2888), .CLK(clk), .Q(\Mem[18][26] ) );
  DFFPOSX1 \Mem_reg[18][25]  ( .D(n2887), .CLK(clk), .Q(\Mem[18][25] ) );
  DFFPOSX1 \Mem_reg[18][24]  ( .D(n2886), .CLK(clk), .Q(\Mem[18][24] ) );
  DFFPOSX1 \Mem_reg[18][23]  ( .D(n2885), .CLK(clk), .Q(\Mem[18][23] ) );
  DFFPOSX1 \Mem_reg[18][22]  ( .D(n2884), .CLK(clk), .Q(\Mem[18][22] ) );
  DFFPOSX1 \Mem_reg[18][21]  ( .D(n2883), .CLK(clk), .Q(\Mem[18][21] ) );
  DFFPOSX1 \Mem_reg[18][20]  ( .D(n2882), .CLK(clk), .Q(\Mem[18][20] ) );
  DFFPOSX1 \Mem_reg[18][19]  ( .D(n2881), .CLK(clk), .Q(\Mem[18][19] ) );
  DFFPOSX1 \Mem_reg[18][18]  ( .D(n2880), .CLK(clk), .Q(\Mem[18][18] ) );
  DFFPOSX1 \Mem_reg[18][17]  ( .D(n2879), .CLK(clk), .Q(\Mem[18][17] ) );
  DFFPOSX1 \Mem_reg[18][16]  ( .D(n2878), .CLK(clk), .Q(\Mem[18][16] ) );
  DFFPOSX1 \Mem_reg[18][15]  ( .D(n2877), .CLK(clk), .Q(\Mem[18][15] ) );
  DFFPOSX1 \Mem_reg[18][14]  ( .D(n2876), .CLK(clk), .Q(\Mem[18][14] ) );
  DFFPOSX1 \Mem_reg[18][13]  ( .D(n2875), .CLK(clk), .Q(\Mem[18][13] ) );
  DFFPOSX1 \Mem_reg[18][12]  ( .D(n2874), .CLK(clk), .Q(\Mem[18][12] ) );
  DFFPOSX1 \Mem_reg[18][11]  ( .D(n2873), .CLK(clk), .Q(\Mem[18][11] ) );
  DFFPOSX1 \Mem_reg[18][10]  ( .D(n2872), .CLK(clk), .Q(\Mem[18][10] ) );
  DFFPOSX1 \Mem_reg[18][9]  ( .D(n2871), .CLK(clk), .Q(\Mem[18][9] ) );
  DFFPOSX1 \Mem_reg[18][8]  ( .D(n2870), .CLK(clk), .Q(\Mem[18][8] ) );
  DFFPOSX1 \Mem_reg[18][7]  ( .D(n2869), .CLK(clk), .Q(\Mem[18][7] ) );
  DFFPOSX1 \Mem_reg[18][6]  ( .D(n2868), .CLK(clk), .Q(\Mem[18][6] ) );
  DFFPOSX1 \Mem_reg[18][5]  ( .D(n2867), .CLK(clk), .Q(\Mem[18][5] ) );
  DFFPOSX1 \Mem_reg[18][4]  ( .D(n2866), .CLK(clk), .Q(\Mem[18][4] ) );
  DFFPOSX1 \Mem_reg[18][3]  ( .D(n2865), .CLK(clk), .Q(\Mem[18][3] ) );
  DFFPOSX1 \Mem_reg[18][2]  ( .D(n2864), .CLK(clk), .Q(\Mem[18][2] ) );
  DFFPOSX1 \Mem_reg[18][1]  ( .D(n2863), .CLK(clk), .Q(\Mem[18][1] ) );
  DFFPOSX1 \Mem_reg[18][0]  ( .D(n2862), .CLK(clk), .Q(\Mem[18][0] ) );
  DFFPOSX1 \Mem_reg[17][31]  ( .D(n2861), .CLK(clk), .Q(\Mem[17][31] ) );
  DFFPOSX1 \Mem_reg[17][30]  ( .D(n2860), .CLK(clk), .Q(\Mem[17][30] ) );
  DFFPOSX1 \Mem_reg[17][29]  ( .D(n2859), .CLK(clk), .Q(\Mem[17][29] ) );
  DFFPOSX1 \Mem_reg[17][28]  ( .D(n2858), .CLK(clk), .Q(\Mem[17][28] ) );
  DFFPOSX1 \Mem_reg[17][27]  ( .D(n2857), .CLK(clk), .Q(\Mem[17][27] ) );
  DFFPOSX1 \Mem_reg[17][26]  ( .D(n2856), .CLK(clk), .Q(\Mem[17][26] ) );
  DFFPOSX1 \Mem_reg[17][25]  ( .D(n2855), .CLK(clk), .Q(\Mem[17][25] ) );
  DFFPOSX1 \Mem_reg[17][24]  ( .D(n2854), .CLK(clk), .Q(\Mem[17][24] ) );
  DFFPOSX1 \Mem_reg[17][23]  ( .D(n2853), .CLK(clk), .Q(\Mem[17][23] ) );
  DFFPOSX1 \Mem_reg[17][22]  ( .D(n2852), .CLK(clk), .Q(\Mem[17][22] ) );
  DFFPOSX1 \Mem_reg[17][21]  ( .D(n2851), .CLK(clk), .Q(\Mem[17][21] ) );
  DFFPOSX1 \Mem_reg[17][20]  ( .D(n2850), .CLK(clk), .Q(\Mem[17][20] ) );
  DFFPOSX1 \Mem_reg[17][19]  ( .D(n2849), .CLK(clk), .Q(\Mem[17][19] ) );
  DFFPOSX1 \Mem_reg[17][18]  ( .D(n2848), .CLK(clk), .Q(\Mem[17][18] ) );
  DFFPOSX1 \Mem_reg[17][17]  ( .D(n2847), .CLK(clk), .Q(\Mem[17][17] ) );
  DFFPOSX1 \Mem_reg[17][16]  ( .D(n2846), .CLK(clk), .Q(\Mem[17][16] ) );
  DFFPOSX1 \Mem_reg[17][15]  ( .D(n2845), .CLK(clk), .Q(\Mem[17][15] ) );
  DFFPOSX1 \Mem_reg[17][14]  ( .D(n2844), .CLK(clk), .Q(\Mem[17][14] ) );
  DFFPOSX1 \Mem_reg[17][13]  ( .D(n2843), .CLK(clk), .Q(\Mem[17][13] ) );
  DFFPOSX1 \Mem_reg[17][12]  ( .D(n2842), .CLK(clk), .Q(\Mem[17][12] ) );
  DFFPOSX1 \Mem_reg[17][11]  ( .D(n2841), .CLK(clk), .Q(\Mem[17][11] ) );
  DFFPOSX1 \Mem_reg[17][10]  ( .D(n2840), .CLK(clk), .Q(\Mem[17][10] ) );
  DFFPOSX1 \Mem_reg[17][9]  ( .D(n2839), .CLK(clk), .Q(\Mem[17][9] ) );
  DFFPOSX1 \Mem_reg[17][8]  ( .D(n2838), .CLK(clk), .Q(\Mem[17][8] ) );
  DFFPOSX1 \Mem_reg[17][7]  ( .D(n2837), .CLK(clk), .Q(\Mem[17][7] ) );
  DFFPOSX1 \Mem_reg[17][6]  ( .D(n2836), .CLK(clk), .Q(\Mem[17][6] ) );
  DFFPOSX1 \Mem_reg[17][5]  ( .D(n2835), .CLK(clk), .Q(\Mem[17][5] ) );
  DFFPOSX1 \Mem_reg[17][4]  ( .D(n2834), .CLK(clk), .Q(\Mem[17][4] ) );
  DFFPOSX1 \Mem_reg[17][3]  ( .D(n2833), .CLK(clk), .Q(\Mem[17][3] ) );
  DFFPOSX1 \Mem_reg[17][2]  ( .D(n2832), .CLK(clk), .Q(\Mem[17][2] ) );
  DFFPOSX1 \Mem_reg[17][1]  ( .D(n2831), .CLK(clk), .Q(\Mem[17][1] ) );
  DFFPOSX1 \Mem_reg[17][0]  ( .D(n2830), .CLK(clk), .Q(\Mem[17][0] ) );
  DFFPOSX1 \Mem_reg[16][31]  ( .D(n2829), .CLK(clk), .Q(\Mem[16][31] ) );
  DFFPOSX1 \Mem_reg[16][30]  ( .D(n2828), .CLK(clk), .Q(\Mem[16][30] ) );
  DFFPOSX1 \Mem_reg[16][29]  ( .D(n2827), .CLK(clk), .Q(\Mem[16][29] ) );
  DFFPOSX1 \Mem_reg[16][28]  ( .D(n2826), .CLK(clk), .Q(\Mem[16][28] ) );
  DFFPOSX1 \Mem_reg[16][27]  ( .D(n2825), .CLK(clk), .Q(\Mem[16][27] ) );
  DFFPOSX1 \Mem_reg[16][26]  ( .D(n2824), .CLK(clk), .Q(\Mem[16][26] ) );
  DFFPOSX1 \Mem_reg[16][25]  ( .D(n2823), .CLK(clk), .Q(\Mem[16][25] ) );
  DFFPOSX1 \Mem_reg[16][24]  ( .D(n2822), .CLK(clk), .Q(\Mem[16][24] ) );
  DFFPOSX1 \Mem_reg[16][23]  ( .D(n2821), .CLK(clk), .Q(\Mem[16][23] ) );
  DFFPOSX1 \Mem_reg[16][22]  ( .D(n2820), .CLK(clk), .Q(\Mem[16][22] ) );
  DFFPOSX1 \Mem_reg[16][21]  ( .D(n2819), .CLK(clk), .Q(\Mem[16][21] ) );
  DFFPOSX1 \Mem_reg[16][20]  ( .D(n2818), .CLK(clk), .Q(\Mem[16][20] ) );
  DFFPOSX1 \Mem_reg[16][19]  ( .D(n2817), .CLK(clk), .Q(\Mem[16][19] ) );
  DFFPOSX1 \Mem_reg[16][18]  ( .D(n2816), .CLK(clk), .Q(\Mem[16][18] ) );
  DFFPOSX1 \Mem_reg[16][17]  ( .D(n2815), .CLK(clk), .Q(\Mem[16][17] ) );
  DFFPOSX1 \Mem_reg[16][16]  ( .D(n2814), .CLK(clk), .Q(\Mem[16][16] ) );
  DFFPOSX1 \Mem_reg[16][15]  ( .D(n2813), .CLK(clk), .Q(\Mem[16][15] ) );
  DFFPOSX1 \Mem_reg[16][14]  ( .D(n2812), .CLK(clk), .Q(\Mem[16][14] ) );
  DFFPOSX1 \Mem_reg[16][13]  ( .D(n2811), .CLK(clk), .Q(\Mem[16][13] ) );
  DFFPOSX1 \Mem_reg[16][12]  ( .D(n2810), .CLK(clk), .Q(\Mem[16][12] ) );
  DFFPOSX1 \Mem_reg[16][11]  ( .D(n2809), .CLK(clk), .Q(\Mem[16][11] ) );
  DFFPOSX1 \Mem_reg[16][10]  ( .D(n2808), .CLK(clk), .Q(\Mem[16][10] ) );
  DFFPOSX1 \Mem_reg[16][9]  ( .D(n2807), .CLK(clk), .Q(\Mem[16][9] ) );
  DFFPOSX1 \Mem_reg[16][8]  ( .D(n2806), .CLK(clk), .Q(\Mem[16][8] ) );
  DFFPOSX1 \Mem_reg[16][7]  ( .D(n2805), .CLK(clk), .Q(\Mem[16][7] ) );
  DFFPOSX1 \Mem_reg[16][6]  ( .D(n2804), .CLK(clk), .Q(\Mem[16][6] ) );
  DFFPOSX1 \Mem_reg[16][5]  ( .D(n2803), .CLK(clk), .Q(\Mem[16][5] ) );
  DFFPOSX1 \Mem_reg[16][4]  ( .D(n2802), .CLK(clk), .Q(\Mem[16][4] ) );
  DFFPOSX1 \Mem_reg[16][3]  ( .D(n2801), .CLK(clk), .Q(\Mem[16][3] ) );
  DFFPOSX1 \Mem_reg[16][2]  ( .D(n2800), .CLK(clk), .Q(\Mem[16][2] ) );
  DFFPOSX1 \Mem_reg[16][1]  ( .D(n2799), .CLK(clk), .Q(\Mem[16][1] ) );
  DFFPOSX1 \Mem_reg[16][0]  ( .D(n2798), .CLK(clk), .Q(\Mem[16][0] ) );
  DFFPOSX1 \Mem_reg[15][31]  ( .D(n2797), .CLK(clk), .Q(\Mem[15][31] ) );
  DFFPOSX1 \Mem_reg[15][30]  ( .D(n2796), .CLK(clk), .Q(\Mem[15][30] ) );
  DFFPOSX1 \Mem_reg[15][29]  ( .D(n2795), .CLK(clk), .Q(\Mem[15][29] ) );
  DFFPOSX1 \Mem_reg[15][28]  ( .D(n2794), .CLK(clk), .Q(\Mem[15][28] ) );
  DFFPOSX1 \Mem_reg[15][27]  ( .D(n2793), .CLK(clk), .Q(\Mem[15][27] ) );
  DFFPOSX1 \Mem_reg[15][26]  ( .D(n2792), .CLK(clk), .Q(\Mem[15][26] ) );
  DFFPOSX1 \Mem_reg[15][25]  ( .D(n2791), .CLK(clk), .Q(\Mem[15][25] ) );
  DFFPOSX1 \Mem_reg[15][24]  ( .D(n2790), .CLK(clk), .Q(\Mem[15][24] ) );
  DFFPOSX1 \Mem_reg[15][23]  ( .D(n2789), .CLK(clk), .Q(\Mem[15][23] ) );
  DFFPOSX1 \Mem_reg[15][22]  ( .D(n2788), .CLK(clk), .Q(\Mem[15][22] ) );
  DFFPOSX1 \Mem_reg[15][21]  ( .D(n2787), .CLK(clk), .Q(\Mem[15][21] ) );
  DFFPOSX1 \Mem_reg[15][20]  ( .D(n2786), .CLK(clk), .Q(\Mem[15][20] ) );
  DFFPOSX1 \Mem_reg[15][19]  ( .D(n2785), .CLK(clk), .Q(\Mem[15][19] ) );
  DFFPOSX1 \Mem_reg[15][18]  ( .D(n2784), .CLK(clk), .Q(\Mem[15][18] ) );
  DFFPOSX1 \Mem_reg[15][17]  ( .D(n2783), .CLK(clk), .Q(\Mem[15][17] ) );
  DFFPOSX1 \Mem_reg[15][16]  ( .D(n2782), .CLK(clk), .Q(\Mem[15][16] ) );
  DFFPOSX1 \Mem_reg[15][15]  ( .D(n2781), .CLK(clk), .Q(\Mem[15][15] ) );
  DFFPOSX1 \Mem_reg[15][14]  ( .D(n2780), .CLK(clk), .Q(\Mem[15][14] ) );
  DFFPOSX1 \Mem_reg[15][13]  ( .D(n2779), .CLK(clk), .Q(\Mem[15][13] ) );
  DFFPOSX1 \Mem_reg[15][12]  ( .D(n2778), .CLK(clk), .Q(\Mem[15][12] ) );
  DFFPOSX1 \Mem_reg[15][11]  ( .D(n2777), .CLK(clk), .Q(\Mem[15][11] ) );
  DFFPOSX1 \Mem_reg[15][10]  ( .D(n2776), .CLK(clk), .Q(\Mem[15][10] ) );
  DFFPOSX1 \Mem_reg[15][9]  ( .D(n2775), .CLK(clk), .Q(\Mem[15][9] ) );
  DFFPOSX1 \Mem_reg[15][8]  ( .D(n2774), .CLK(clk), .Q(\Mem[15][8] ) );
  DFFPOSX1 \Mem_reg[15][7]  ( .D(n2773), .CLK(clk), .Q(\Mem[15][7] ) );
  DFFPOSX1 \Mem_reg[15][6]  ( .D(n2772), .CLK(clk), .Q(\Mem[15][6] ) );
  DFFPOSX1 \Mem_reg[15][5]  ( .D(n2771), .CLK(clk), .Q(\Mem[15][5] ) );
  DFFPOSX1 \Mem_reg[15][4]  ( .D(n2770), .CLK(clk), .Q(\Mem[15][4] ) );
  DFFPOSX1 \Mem_reg[15][3]  ( .D(n2769), .CLK(clk), .Q(\Mem[15][3] ) );
  DFFPOSX1 \Mem_reg[15][2]  ( .D(n2768), .CLK(clk), .Q(\Mem[15][2] ) );
  DFFPOSX1 \Mem_reg[15][1]  ( .D(n2767), .CLK(clk), .Q(\Mem[15][1] ) );
  DFFPOSX1 \Mem_reg[15][0]  ( .D(n2766), .CLK(clk), .Q(\Mem[15][0] ) );
  DFFPOSX1 \Mem_reg[14][31]  ( .D(n2765), .CLK(clk), .Q(\Mem[14][31] ) );
  DFFPOSX1 \Mem_reg[14][30]  ( .D(n2764), .CLK(clk), .Q(\Mem[14][30] ) );
  DFFPOSX1 \Mem_reg[14][29]  ( .D(n2763), .CLK(clk), .Q(\Mem[14][29] ) );
  DFFPOSX1 \Mem_reg[14][28]  ( .D(n2762), .CLK(clk), .Q(\Mem[14][28] ) );
  DFFPOSX1 \Mem_reg[14][27]  ( .D(n2761), .CLK(clk), .Q(\Mem[14][27] ) );
  DFFPOSX1 \Mem_reg[14][26]  ( .D(n2760), .CLK(clk), .Q(\Mem[14][26] ) );
  DFFPOSX1 \Mem_reg[14][25]  ( .D(n2759), .CLK(clk), .Q(\Mem[14][25] ) );
  DFFPOSX1 \Mem_reg[14][24]  ( .D(n2758), .CLK(clk), .Q(\Mem[14][24] ) );
  DFFPOSX1 \Mem_reg[14][23]  ( .D(n2757), .CLK(clk), .Q(\Mem[14][23] ) );
  DFFPOSX1 \Mem_reg[14][22]  ( .D(n2756), .CLK(clk), .Q(\Mem[14][22] ) );
  DFFPOSX1 \Mem_reg[14][21]  ( .D(n2755), .CLK(clk), .Q(\Mem[14][21] ) );
  DFFPOSX1 \Mem_reg[14][20]  ( .D(n2754), .CLK(clk), .Q(\Mem[14][20] ) );
  DFFPOSX1 \Mem_reg[14][19]  ( .D(n2753), .CLK(clk), .Q(\Mem[14][19] ) );
  DFFPOSX1 \Mem_reg[14][18]  ( .D(n2752), .CLK(clk), .Q(\Mem[14][18] ) );
  DFFPOSX1 \Mem_reg[14][17]  ( .D(n2751), .CLK(clk), .Q(\Mem[14][17] ) );
  DFFPOSX1 \Mem_reg[14][16]  ( .D(n2750), .CLK(clk), .Q(\Mem[14][16] ) );
  DFFPOSX1 \Mem_reg[14][15]  ( .D(n2749), .CLK(clk), .Q(\Mem[14][15] ) );
  DFFPOSX1 \Mem_reg[14][14]  ( .D(n2748), .CLK(clk), .Q(\Mem[14][14] ) );
  DFFPOSX1 \Mem_reg[14][13]  ( .D(n2747), .CLK(clk), .Q(\Mem[14][13] ) );
  DFFPOSX1 \Mem_reg[14][12]  ( .D(n2746), .CLK(clk), .Q(\Mem[14][12] ) );
  DFFPOSX1 \Mem_reg[14][11]  ( .D(n2745), .CLK(clk), .Q(\Mem[14][11] ) );
  DFFPOSX1 \Mem_reg[14][10]  ( .D(n2744), .CLK(clk), .Q(\Mem[14][10] ) );
  DFFPOSX1 \Mem_reg[14][9]  ( .D(n2743), .CLK(clk), .Q(\Mem[14][9] ) );
  DFFPOSX1 \Mem_reg[14][8]  ( .D(n2742), .CLK(clk), .Q(\Mem[14][8] ) );
  DFFPOSX1 \Mem_reg[14][7]  ( .D(n2741), .CLK(clk), .Q(\Mem[14][7] ) );
  DFFPOSX1 \Mem_reg[14][6]  ( .D(n2740), .CLK(clk), .Q(\Mem[14][6] ) );
  DFFPOSX1 \Mem_reg[14][5]  ( .D(n2739), .CLK(clk), .Q(\Mem[14][5] ) );
  DFFPOSX1 \Mem_reg[14][4]  ( .D(n2738), .CLK(clk), .Q(\Mem[14][4] ) );
  DFFPOSX1 \Mem_reg[14][3]  ( .D(n2737), .CLK(clk), .Q(\Mem[14][3] ) );
  DFFPOSX1 \Mem_reg[14][2]  ( .D(n2736), .CLK(clk), .Q(\Mem[14][2] ) );
  DFFPOSX1 \Mem_reg[14][1]  ( .D(n2735), .CLK(clk), .Q(\Mem[14][1] ) );
  DFFPOSX1 \Mem_reg[14][0]  ( .D(n2734), .CLK(clk), .Q(\Mem[14][0] ) );
  DFFPOSX1 \Mem_reg[13][31]  ( .D(n2733), .CLK(clk), .Q(\Mem[13][31] ) );
  DFFPOSX1 \Mem_reg[13][30]  ( .D(n2732), .CLK(clk), .Q(\Mem[13][30] ) );
  DFFPOSX1 \Mem_reg[13][29]  ( .D(n2731), .CLK(clk), .Q(\Mem[13][29] ) );
  DFFPOSX1 \Mem_reg[13][28]  ( .D(n2730), .CLK(clk), .Q(\Mem[13][28] ) );
  DFFPOSX1 \Mem_reg[13][27]  ( .D(n2729), .CLK(clk), .Q(\Mem[13][27] ) );
  DFFPOSX1 \Mem_reg[13][26]  ( .D(n2728), .CLK(clk), .Q(\Mem[13][26] ) );
  DFFPOSX1 \Mem_reg[13][25]  ( .D(n2727), .CLK(clk), .Q(\Mem[13][25] ) );
  DFFPOSX1 \Mem_reg[13][24]  ( .D(n2726), .CLK(clk), .Q(\Mem[13][24] ) );
  DFFPOSX1 \Mem_reg[13][23]  ( .D(n2725), .CLK(clk), .Q(\Mem[13][23] ) );
  DFFPOSX1 \Mem_reg[13][22]  ( .D(n2724), .CLK(clk), .Q(\Mem[13][22] ) );
  DFFPOSX1 \Mem_reg[13][21]  ( .D(n2723), .CLK(clk), .Q(\Mem[13][21] ) );
  DFFPOSX1 \Mem_reg[13][20]  ( .D(n2722), .CLK(clk), .Q(\Mem[13][20] ) );
  DFFPOSX1 \Mem_reg[13][19]  ( .D(n2721), .CLK(clk), .Q(\Mem[13][19] ) );
  DFFPOSX1 \Mem_reg[13][18]  ( .D(n2720), .CLK(clk), .Q(\Mem[13][18] ) );
  DFFPOSX1 \Mem_reg[13][17]  ( .D(n2719), .CLK(clk), .Q(\Mem[13][17] ) );
  DFFPOSX1 \Mem_reg[13][16]  ( .D(n2718), .CLK(clk), .Q(\Mem[13][16] ) );
  DFFPOSX1 \Mem_reg[13][15]  ( .D(n2717), .CLK(clk), .Q(\Mem[13][15] ) );
  DFFPOSX1 \Mem_reg[13][14]  ( .D(n2716), .CLK(clk), .Q(\Mem[13][14] ) );
  DFFPOSX1 \Mem_reg[13][13]  ( .D(n2715), .CLK(clk), .Q(\Mem[13][13] ) );
  DFFPOSX1 \Mem_reg[13][12]  ( .D(n2714), .CLK(clk), .Q(\Mem[13][12] ) );
  DFFPOSX1 \Mem_reg[13][11]  ( .D(n2713), .CLK(clk), .Q(\Mem[13][11] ) );
  DFFPOSX1 \Mem_reg[13][10]  ( .D(n2712), .CLK(clk), .Q(\Mem[13][10] ) );
  DFFPOSX1 \Mem_reg[13][9]  ( .D(n2711), .CLK(clk), .Q(\Mem[13][9] ) );
  DFFPOSX1 \Mem_reg[13][8]  ( .D(n2710), .CLK(clk), .Q(\Mem[13][8] ) );
  DFFPOSX1 \Mem_reg[13][7]  ( .D(n2709), .CLK(clk), .Q(\Mem[13][7] ) );
  DFFPOSX1 \Mem_reg[13][6]  ( .D(n2708), .CLK(clk), .Q(\Mem[13][6] ) );
  DFFPOSX1 \Mem_reg[13][5]  ( .D(n2707), .CLK(clk), .Q(\Mem[13][5] ) );
  DFFPOSX1 \Mem_reg[13][4]  ( .D(n2706), .CLK(clk), .Q(\Mem[13][4] ) );
  DFFPOSX1 \Mem_reg[13][3]  ( .D(n2705), .CLK(clk), .Q(\Mem[13][3] ) );
  DFFPOSX1 \Mem_reg[13][2]  ( .D(n2704), .CLK(clk), .Q(\Mem[13][2] ) );
  DFFPOSX1 \Mem_reg[13][1]  ( .D(n2703), .CLK(clk), .Q(\Mem[13][1] ) );
  DFFPOSX1 \Mem_reg[13][0]  ( .D(n2702), .CLK(clk), .Q(\Mem[13][0] ) );
  DFFPOSX1 \Mem_reg[12][31]  ( .D(n2701), .CLK(clk), .Q(\Mem[12][31] ) );
  DFFPOSX1 \Mem_reg[12][30]  ( .D(n2700), .CLK(clk), .Q(\Mem[12][30] ) );
  DFFPOSX1 \Mem_reg[12][29]  ( .D(n2699), .CLK(clk), .Q(\Mem[12][29] ) );
  DFFPOSX1 \Mem_reg[12][28]  ( .D(n2698), .CLK(clk), .Q(\Mem[12][28] ) );
  DFFPOSX1 \Mem_reg[12][27]  ( .D(n2697), .CLK(clk), .Q(\Mem[12][27] ) );
  DFFPOSX1 \Mem_reg[12][26]  ( .D(n2696), .CLK(clk), .Q(\Mem[12][26] ) );
  DFFPOSX1 \Mem_reg[12][25]  ( .D(n2695), .CLK(clk), .Q(\Mem[12][25] ) );
  DFFPOSX1 \Mem_reg[12][24]  ( .D(n2694), .CLK(clk), .Q(\Mem[12][24] ) );
  DFFPOSX1 \Mem_reg[12][23]  ( .D(n2693), .CLK(clk), .Q(\Mem[12][23] ) );
  DFFPOSX1 \Mem_reg[12][22]  ( .D(n2692), .CLK(clk), .Q(\Mem[12][22] ) );
  DFFPOSX1 \Mem_reg[12][21]  ( .D(n2691), .CLK(clk), .Q(\Mem[12][21] ) );
  DFFPOSX1 \Mem_reg[12][20]  ( .D(n2690), .CLK(clk), .Q(\Mem[12][20] ) );
  DFFPOSX1 \Mem_reg[12][19]  ( .D(n2689), .CLK(clk), .Q(\Mem[12][19] ) );
  DFFPOSX1 \Mem_reg[12][18]  ( .D(n2688), .CLK(clk), .Q(\Mem[12][18] ) );
  DFFPOSX1 \Mem_reg[12][17]  ( .D(n2687), .CLK(clk), .Q(\Mem[12][17] ) );
  DFFPOSX1 \Mem_reg[12][16]  ( .D(n2686), .CLK(clk), .Q(\Mem[12][16] ) );
  DFFPOSX1 \Mem_reg[12][15]  ( .D(n2685), .CLK(clk), .Q(\Mem[12][15] ) );
  DFFPOSX1 \Mem_reg[12][14]  ( .D(n2684), .CLK(clk), .Q(\Mem[12][14] ) );
  DFFPOSX1 \Mem_reg[12][13]  ( .D(n2683), .CLK(clk), .Q(\Mem[12][13] ) );
  DFFPOSX1 \Mem_reg[12][12]  ( .D(n2682), .CLK(clk), .Q(\Mem[12][12] ) );
  DFFPOSX1 \Mem_reg[12][11]  ( .D(n2681), .CLK(clk), .Q(\Mem[12][11] ) );
  DFFPOSX1 \Mem_reg[12][10]  ( .D(n2680), .CLK(clk), .Q(\Mem[12][10] ) );
  DFFPOSX1 \Mem_reg[12][9]  ( .D(n2679), .CLK(clk), .Q(\Mem[12][9] ) );
  DFFPOSX1 \Mem_reg[12][8]  ( .D(n2678), .CLK(clk), .Q(\Mem[12][8] ) );
  DFFPOSX1 \Mem_reg[12][7]  ( .D(n2677), .CLK(clk), .Q(\Mem[12][7] ) );
  DFFPOSX1 \Mem_reg[12][6]  ( .D(n2676), .CLK(clk), .Q(\Mem[12][6] ) );
  DFFPOSX1 \Mem_reg[12][5]  ( .D(n2675), .CLK(clk), .Q(\Mem[12][5] ) );
  DFFPOSX1 \Mem_reg[12][4]  ( .D(n2674), .CLK(clk), .Q(\Mem[12][4] ) );
  DFFPOSX1 \Mem_reg[12][3]  ( .D(n2673), .CLK(clk), .Q(\Mem[12][3] ) );
  DFFPOSX1 \Mem_reg[12][2]  ( .D(n2672), .CLK(clk), .Q(\Mem[12][2] ) );
  DFFPOSX1 \Mem_reg[12][1]  ( .D(n2671), .CLK(clk), .Q(\Mem[12][1] ) );
  DFFPOSX1 \Mem_reg[12][0]  ( .D(n2670), .CLK(clk), .Q(\Mem[12][0] ) );
  DFFPOSX1 \Mem_reg[11][31]  ( .D(n2669), .CLK(clk), .Q(\Mem[11][31] ) );
  DFFPOSX1 \Mem_reg[11][30]  ( .D(n2668), .CLK(clk), .Q(\Mem[11][30] ) );
  DFFPOSX1 \Mem_reg[11][29]  ( .D(n2667), .CLK(clk), .Q(\Mem[11][29] ) );
  DFFPOSX1 \Mem_reg[11][28]  ( .D(n2666), .CLK(clk), .Q(\Mem[11][28] ) );
  DFFPOSX1 \Mem_reg[11][27]  ( .D(n2665), .CLK(clk), .Q(\Mem[11][27] ) );
  DFFPOSX1 \Mem_reg[11][26]  ( .D(n2664), .CLK(clk), .Q(\Mem[11][26] ) );
  DFFPOSX1 \Mem_reg[11][25]  ( .D(n2663), .CLK(clk), .Q(\Mem[11][25] ) );
  DFFPOSX1 \Mem_reg[11][24]  ( .D(n2662), .CLK(clk), .Q(\Mem[11][24] ) );
  DFFPOSX1 \Mem_reg[11][23]  ( .D(n2661), .CLK(clk), .Q(\Mem[11][23] ) );
  DFFPOSX1 \Mem_reg[11][22]  ( .D(n2660), .CLK(clk), .Q(\Mem[11][22] ) );
  DFFPOSX1 \Mem_reg[11][21]  ( .D(n2659), .CLK(clk), .Q(\Mem[11][21] ) );
  DFFPOSX1 \Mem_reg[11][20]  ( .D(n2658), .CLK(clk), .Q(\Mem[11][20] ) );
  DFFPOSX1 \Mem_reg[11][19]  ( .D(n2657), .CLK(clk), .Q(\Mem[11][19] ) );
  DFFPOSX1 \Mem_reg[11][18]  ( .D(n2656), .CLK(clk), .Q(\Mem[11][18] ) );
  DFFPOSX1 \Mem_reg[11][17]  ( .D(n2655), .CLK(clk), .Q(\Mem[11][17] ) );
  DFFPOSX1 \Mem_reg[11][16]  ( .D(n2654), .CLK(clk), .Q(\Mem[11][16] ) );
  DFFPOSX1 \Mem_reg[11][15]  ( .D(n2653), .CLK(clk), .Q(\Mem[11][15] ) );
  DFFPOSX1 \Mem_reg[11][14]  ( .D(n2652), .CLK(clk), .Q(\Mem[11][14] ) );
  DFFPOSX1 \Mem_reg[11][13]  ( .D(n2651), .CLK(clk), .Q(\Mem[11][13] ) );
  DFFPOSX1 \Mem_reg[11][12]  ( .D(n2650), .CLK(clk), .Q(\Mem[11][12] ) );
  DFFPOSX1 \Mem_reg[11][11]  ( .D(n2649), .CLK(clk), .Q(\Mem[11][11] ) );
  DFFPOSX1 \Mem_reg[11][10]  ( .D(n2648), .CLK(clk), .Q(\Mem[11][10] ) );
  DFFPOSX1 \Mem_reg[11][9]  ( .D(n2647), .CLK(clk), .Q(\Mem[11][9] ) );
  DFFPOSX1 \Mem_reg[11][8]  ( .D(n2646), .CLK(clk), .Q(\Mem[11][8] ) );
  DFFPOSX1 \Mem_reg[11][7]  ( .D(n2645), .CLK(clk), .Q(\Mem[11][7] ) );
  DFFPOSX1 \Mem_reg[11][6]  ( .D(n2644), .CLK(clk), .Q(\Mem[11][6] ) );
  DFFPOSX1 \Mem_reg[11][5]  ( .D(n2643), .CLK(clk), .Q(\Mem[11][5] ) );
  DFFPOSX1 \Mem_reg[11][4]  ( .D(n2642), .CLK(clk), .Q(\Mem[11][4] ) );
  DFFPOSX1 \Mem_reg[11][3]  ( .D(n2641), .CLK(clk), .Q(\Mem[11][3] ) );
  DFFPOSX1 \Mem_reg[11][2]  ( .D(n2640), .CLK(clk), .Q(\Mem[11][2] ) );
  DFFPOSX1 \Mem_reg[11][1]  ( .D(n2639), .CLK(clk), .Q(\Mem[11][1] ) );
  DFFPOSX1 \Mem_reg[11][0]  ( .D(n2638), .CLK(clk), .Q(\Mem[11][0] ) );
  DFFPOSX1 \Mem_reg[10][31]  ( .D(n2637), .CLK(clk), .Q(\Mem[10][31] ) );
  DFFPOSX1 \Mem_reg[10][30]  ( .D(n2636), .CLK(clk), .Q(\Mem[10][30] ) );
  DFFPOSX1 \Mem_reg[10][29]  ( .D(n2635), .CLK(clk), .Q(\Mem[10][29] ) );
  DFFPOSX1 \Mem_reg[10][28]  ( .D(n2634), .CLK(clk), .Q(\Mem[10][28] ) );
  DFFPOSX1 \Mem_reg[10][27]  ( .D(n2633), .CLK(clk), .Q(\Mem[10][27] ) );
  DFFPOSX1 \Mem_reg[10][26]  ( .D(n2632), .CLK(clk), .Q(\Mem[10][26] ) );
  DFFPOSX1 \Mem_reg[10][25]  ( .D(n2631), .CLK(clk), .Q(\Mem[10][25] ) );
  DFFPOSX1 \Mem_reg[10][24]  ( .D(n2630), .CLK(clk), .Q(\Mem[10][24] ) );
  DFFPOSX1 \Mem_reg[10][23]  ( .D(n2629), .CLK(clk), .Q(\Mem[10][23] ) );
  DFFPOSX1 \Mem_reg[10][22]  ( .D(n2628), .CLK(clk), .Q(\Mem[10][22] ) );
  DFFPOSX1 \Mem_reg[10][21]  ( .D(n2627), .CLK(clk), .Q(\Mem[10][21] ) );
  DFFPOSX1 \Mem_reg[10][20]  ( .D(n2626), .CLK(clk), .Q(\Mem[10][20] ) );
  DFFPOSX1 \Mem_reg[10][19]  ( .D(n2625), .CLK(clk), .Q(\Mem[10][19] ) );
  DFFPOSX1 \Mem_reg[10][18]  ( .D(n2624), .CLK(clk), .Q(\Mem[10][18] ) );
  DFFPOSX1 \Mem_reg[10][17]  ( .D(n2623), .CLK(clk), .Q(\Mem[10][17] ) );
  DFFPOSX1 \Mem_reg[10][16]  ( .D(n2622), .CLK(clk), .Q(\Mem[10][16] ) );
  DFFPOSX1 \Mem_reg[10][15]  ( .D(n2621), .CLK(clk), .Q(\Mem[10][15] ) );
  DFFPOSX1 \Mem_reg[10][14]  ( .D(n2620), .CLK(clk), .Q(\Mem[10][14] ) );
  DFFPOSX1 \Mem_reg[10][13]  ( .D(n2619), .CLK(clk), .Q(\Mem[10][13] ) );
  DFFPOSX1 \Mem_reg[10][12]  ( .D(n2618), .CLK(clk), .Q(\Mem[10][12] ) );
  DFFPOSX1 \Mem_reg[10][11]  ( .D(n2617), .CLK(clk), .Q(\Mem[10][11] ) );
  DFFPOSX1 \Mem_reg[10][10]  ( .D(n2616), .CLK(clk), .Q(\Mem[10][10] ) );
  DFFPOSX1 \Mem_reg[10][9]  ( .D(n2615), .CLK(clk), .Q(\Mem[10][9] ) );
  DFFPOSX1 \Mem_reg[10][8]  ( .D(n2614), .CLK(clk), .Q(\Mem[10][8] ) );
  DFFPOSX1 \Mem_reg[10][7]  ( .D(n2613), .CLK(clk), .Q(\Mem[10][7] ) );
  DFFPOSX1 \Mem_reg[10][6]  ( .D(n2612), .CLK(clk), .Q(\Mem[10][6] ) );
  DFFPOSX1 \Mem_reg[10][5]  ( .D(n2611), .CLK(clk), .Q(\Mem[10][5] ) );
  DFFPOSX1 \Mem_reg[10][4]  ( .D(n2610), .CLK(clk), .Q(\Mem[10][4] ) );
  DFFPOSX1 \Mem_reg[10][3]  ( .D(n2609), .CLK(clk), .Q(\Mem[10][3] ) );
  DFFPOSX1 \Mem_reg[10][2]  ( .D(n2608), .CLK(clk), .Q(\Mem[10][2] ) );
  DFFPOSX1 \Mem_reg[10][1]  ( .D(n2607), .CLK(clk), .Q(\Mem[10][1] ) );
  DFFPOSX1 \Mem_reg[10][0]  ( .D(n2606), .CLK(clk), .Q(\Mem[10][0] ) );
  DFFPOSX1 \Mem_reg[9][31]  ( .D(n2605), .CLK(clk), .Q(\Mem[9][31] ) );
  DFFPOSX1 \Mem_reg[9][30]  ( .D(n2604), .CLK(clk), .Q(\Mem[9][30] ) );
  DFFPOSX1 \Mem_reg[9][29]  ( .D(n2603), .CLK(clk), .Q(\Mem[9][29] ) );
  DFFPOSX1 \Mem_reg[9][28]  ( .D(n2602), .CLK(clk), .Q(\Mem[9][28] ) );
  DFFPOSX1 \Mem_reg[9][27]  ( .D(n2601), .CLK(clk), .Q(\Mem[9][27] ) );
  DFFPOSX1 \Mem_reg[9][26]  ( .D(n2600), .CLK(clk), .Q(\Mem[9][26] ) );
  DFFPOSX1 \Mem_reg[9][25]  ( .D(n2599), .CLK(clk), .Q(\Mem[9][25] ) );
  DFFPOSX1 \Mem_reg[9][24]  ( .D(n2598), .CLK(clk), .Q(\Mem[9][24] ) );
  DFFPOSX1 \Mem_reg[9][23]  ( .D(n2597), .CLK(clk), .Q(\Mem[9][23] ) );
  DFFPOSX1 \Mem_reg[9][22]  ( .D(n2596), .CLK(clk), .Q(\Mem[9][22] ) );
  DFFPOSX1 \Mem_reg[9][21]  ( .D(n2595), .CLK(clk), .Q(\Mem[9][21] ) );
  DFFPOSX1 \Mem_reg[9][20]  ( .D(n2594), .CLK(clk), .Q(\Mem[9][20] ) );
  DFFPOSX1 \Mem_reg[9][19]  ( .D(n2593), .CLK(clk), .Q(\Mem[9][19] ) );
  DFFPOSX1 \Mem_reg[9][18]  ( .D(n2592), .CLK(clk), .Q(\Mem[9][18] ) );
  DFFPOSX1 \Mem_reg[9][17]  ( .D(n2591), .CLK(clk), .Q(\Mem[9][17] ) );
  DFFPOSX1 \Mem_reg[9][16]  ( .D(n2590), .CLK(clk), .Q(\Mem[9][16] ) );
  DFFPOSX1 \Mem_reg[9][15]  ( .D(n2589), .CLK(clk), .Q(\Mem[9][15] ) );
  DFFPOSX1 \Mem_reg[9][14]  ( .D(n2588), .CLK(clk), .Q(\Mem[9][14] ) );
  DFFPOSX1 \Mem_reg[9][13]  ( .D(n2587), .CLK(clk), .Q(\Mem[9][13] ) );
  DFFPOSX1 \Mem_reg[9][12]  ( .D(n2586), .CLK(clk), .Q(\Mem[9][12] ) );
  DFFPOSX1 \Mem_reg[9][11]  ( .D(n2585), .CLK(clk), .Q(\Mem[9][11] ) );
  DFFPOSX1 \Mem_reg[9][10]  ( .D(n2584), .CLK(clk), .Q(\Mem[9][10] ) );
  DFFPOSX1 \Mem_reg[9][9]  ( .D(n2583), .CLK(clk), .Q(\Mem[9][9] ) );
  DFFPOSX1 \Mem_reg[9][8]  ( .D(n2582), .CLK(clk), .Q(\Mem[9][8] ) );
  DFFPOSX1 \Mem_reg[9][7]  ( .D(n2581), .CLK(clk), .Q(\Mem[9][7] ) );
  DFFPOSX1 \Mem_reg[9][6]  ( .D(n2580), .CLK(clk), .Q(\Mem[9][6] ) );
  DFFPOSX1 \Mem_reg[9][5]  ( .D(n2579), .CLK(clk), .Q(\Mem[9][5] ) );
  DFFPOSX1 \Mem_reg[9][4]  ( .D(n2578), .CLK(clk), .Q(\Mem[9][4] ) );
  DFFPOSX1 \Mem_reg[9][3]  ( .D(n2577), .CLK(clk), .Q(\Mem[9][3] ) );
  DFFPOSX1 \Mem_reg[9][2]  ( .D(n2576), .CLK(clk), .Q(\Mem[9][2] ) );
  DFFPOSX1 \Mem_reg[9][1]  ( .D(n2575), .CLK(clk), .Q(\Mem[9][1] ) );
  DFFPOSX1 \Mem_reg[9][0]  ( .D(n2574), .CLK(clk), .Q(\Mem[9][0] ) );
  DFFPOSX1 \Mem_reg[8][31]  ( .D(n2573), .CLK(clk), .Q(\Mem[8][31] ) );
  DFFPOSX1 \Mem_reg[8][30]  ( .D(n2572), .CLK(clk), .Q(\Mem[8][30] ) );
  DFFPOSX1 \Mem_reg[8][29]  ( .D(n2571), .CLK(clk), .Q(\Mem[8][29] ) );
  DFFPOSX1 \Mem_reg[8][28]  ( .D(n2570), .CLK(clk), .Q(\Mem[8][28] ) );
  DFFPOSX1 \Mem_reg[8][27]  ( .D(n2569), .CLK(clk), .Q(\Mem[8][27] ) );
  DFFPOSX1 \Mem_reg[8][26]  ( .D(n2568), .CLK(clk), .Q(\Mem[8][26] ) );
  DFFPOSX1 \Mem_reg[8][25]  ( .D(n2567), .CLK(clk), .Q(\Mem[8][25] ) );
  DFFPOSX1 \Mem_reg[8][24]  ( .D(n2566), .CLK(clk), .Q(\Mem[8][24] ) );
  DFFPOSX1 \Mem_reg[8][23]  ( .D(n2565), .CLK(clk), .Q(\Mem[8][23] ) );
  DFFPOSX1 \Mem_reg[8][22]  ( .D(n2564), .CLK(clk), .Q(\Mem[8][22] ) );
  DFFPOSX1 \Mem_reg[8][21]  ( .D(n2563), .CLK(clk), .Q(\Mem[8][21] ) );
  DFFPOSX1 \Mem_reg[8][20]  ( .D(n2562), .CLK(clk), .Q(\Mem[8][20] ) );
  DFFPOSX1 \Mem_reg[8][19]  ( .D(n2561), .CLK(clk), .Q(\Mem[8][19] ) );
  DFFPOSX1 \Mem_reg[8][18]  ( .D(n2560), .CLK(clk), .Q(\Mem[8][18] ) );
  DFFPOSX1 \Mem_reg[8][17]  ( .D(n2559), .CLK(clk), .Q(\Mem[8][17] ) );
  DFFPOSX1 \Mem_reg[8][16]  ( .D(n2558), .CLK(clk), .Q(\Mem[8][16] ) );
  DFFPOSX1 \Mem_reg[8][15]  ( .D(n2557), .CLK(clk), .Q(\Mem[8][15] ) );
  DFFPOSX1 \Mem_reg[8][14]  ( .D(n2556), .CLK(clk), .Q(\Mem[8][14] ) );
  DFFPOSX1 \Mem_reg[8][13]  ( .D(n2555), .CLK(clk), .Q(\Mem[8][13] ) );
  DFFPOSX1 \Mem_reg[8][12]  ( .D(n2554), .CLK(clk), .Q(\Mem[8][12] ) );
  DFFPOSX1 \Mem_reg[8][11]  ( .D(n2553), .CLK(clk), .Q(\Mem[8][11] ) );
  DFFPOSX1 \Mem_reg[8][10]  ( .D(n2552), .CLK(clk), .Q(\Mem[8][10] ) );
  DFFPOSX1 \Mem_reg[8][9]  ( .D(n2551), .CLK(clk), .Q(\Mem[8][9] ) );
  DFFPOSX1 \Mem_reg[8][8]  ( .D(n2550), .CLK(clk), .Q(\Mem[8][8] ) );
  DFFPOSX1 \Mem_reg[8][7]  ( .D(n2549), .CLK(clk), .Q(\Mem[8][7] ) );
  DFFPOSX1 \Mem_reg[8][6]  ( .D(n2548), .CLK(clk), .Q(\Mem[8][6] ) );
  DFFPOSX1 \Mem_reg[8][5]  ( .D(n2547), .CLK(clk), .Q(\Mem[8][5] ) );
  DFFPOSX1 \Mem_reg[8][4]  ( .D(n2546), .CLK(clk), .Q(\Mem[8][4] ) );
  DFFPOSX1 \Mem_reg[8][3]  ( .D(n2545), .CLK(clk), .Q(\Mem[8][3] ) );
  DFFPOSX1 \Mem_reg[8][2]  ( .D(n2544), .CLK(clk), .Q(\Mem[8][2] ) );
  DFFPOSX1 \Mem_reg[8][1]  ( .D(n2543), .CLK(clk), .Q(\Mem[8][1] ) );
  DFFPOSX1 \Mem_reg[8][0]  ( .D(n2542), .CLK(clk), .Q(\Mem[8][0] ) );
  DFFPOSX1 \Mem_reg[7][31]  ( .D(n2541), .CLK(clk), .Q(\Mem[7][31] ) );
  DFFPOSX1 \Mem_reg[7][30]  ( .D(n2540), .CLK(clk), .Q(\Mem[7][30] ) );
  DFFPOSX1 \Mem_reg[7][29]  ( .D(n2539), .CLK(clk), .Q(\Mem[7][29] ) );
  DFFPOSX1 \Mem_reg[7][28]  ( .D(n2538), .CLK(clk), .Q(\Mem[7][28] ) );
  DFFPOSX1 \Mem_reg[7][27]  ( .D(n2537), .CLK(clk), .Q(\Mem[7][27] ) );
  DFFPOSX1 \Mem_reg[7][26]  ( .D(n2536), .CLK(clk), .Q(\Mem[7][26] ) );
  DFFPOSX1 \Mem_reg[7][25]  ( .D(n2535), .CLK(clk), .Q(\Mem[7][25] ) );
  DFFPOSX1 \Mem_reg[7][24]  ( .D(n2534), .CLK(clk), .Q(\Mem[7][24] ) );
  DFFPOSX1 \Mem_reg[7][23]  ( .D(n2533), .CLK(clk), .Q(\Mem[7][23] ) );
  DFFPOSX1 \Mem_reg[7][22]  ( .D(n2532), .CLK(clk), .Q(\Mem[7][22] ) );
  DFFPOSX1 \Mem_reg[7][21]  ( .D(n2531), .CLK(clk), .Q(\Mem[7][21] ) );
  DFFPOSX1 \Mem_reg[7][20]  ( .D(n2530), .CLK(clk), .Q(\Mem[7][20] ) );
  DFFPOSX1 \Mem_reg[7][19]  ( .D(n2529), .CLK(clk), .Q(\Mem[7][19] ) );
  DFFPOSX1 \Mem_reg[7][18]  ( .D(n2528), .CLK(clk), .Q(\Mem[7][18] ) );
  DFFPOSX1 \Mem_reg[7][17]  ( .D(n2527), .CLK(clk), .Q(\Mem[7][17] ) );
  DFFPOSX1 \Mem_reg[7][16]  ( .D(n2526), .CLK(clk), .Q(\Mem[7][16] ) );
  DFFPOSX1 \Mem_reg[7][15]  ( .D(n2525), .CLK(clk), .Q(\Mem[7][15] ) );
  DFFPOSX1 \Mem_reg[7][14]  ( .D(n2524), .CLK(clk), .Q(\Mem[7][14] ) );
  DFFPOSX1 \Mem_reg[7][13]  ( .D(n2523), .CLK(clk), .Q(\Mem[7][13] ) );
  DFFPOSX1 \Mem_reg[7][12]  ( .D(n2522), .CLK(clk), .Q(\Mem[7][12] ) );
  DFFPOSX1 \Mem_reg[7][11]  ( .D(n2521), .CLK(clk), .Q(\Mem[7][11] ) );
  DFFPOSX1 \Mem_reg[7][10]  ( .D(n2520), .CLK(clk), .Q(\Mem[7][10] ) );
  DFFPOSX1 \Mem_reg[7][9]  ( .D(n2519), .CLK(clk), .Q(\Mem[7][9] ) );
  DFFPOSX1 \Mem_reg[7][8]  ( .D(n2518), .CLK(clk), .Q(\Mem[7][8] ) );
  DFFPOSX1 \Mem_reg[7][7]  ( .D(n2517), .CLK(clk), .Q(\Mem[7][7] ) );
  DFFPOSX1 \Mem_reg[7][6]  ( .D(n2516), .CLK(clk), .Q(\Mem[7][6] ) );
  DFFPOSX1 \Mem_reg[7][5]  ( .D(n2515), .CLK(clk), .Q(\Mem[7][5] ) );
  DFFPOSX1 \Mem_reg[7][4]  ( .D(n2514), .CLK(clk), .Q(\Mem[7][4] ) );
  DFFPOSX1 \Mem_reg[7][3]  ( .D(n2513), .CLK(clk), .Q(\Mem[7][3] ) );
  DFFPOSX1 \Mem_reg[7][2]  ( .D(n2512), .CLK(clk), .Q(\Mem[7][2] ) );
  DFFPOSX1 \Mem_reg[7][1]  ( .D(n2511), .CLK(clk), .Q(\Mem[7][1] ) );
  DFFPOSX1 \Mem_reg[7][0]  ( .D(n2510), .CLK(clk), .Q(\Mem[7][0] ) );
  DFFPOSX1 \Mem_reg[6][31]  ( .D(n2509), .CLK(clk), .Q(\Mem[6][31] ) );
  DFFPOSX1 \Mem_reg[6][30]  ( .D(n2508), .CLK(clk), .Q(\Mem[6][30] ) );
  DFFPOSX1 \Mem_reg[6][29]  ( .D(n2507), .CLK(clk), .Q(\Mem[6][29] ) );
  DFFPOSX1 \Mem_reg[6][28]  ( .D(n2506), .CLK(clk), .Q(\Mem[6][28] ) );
  DFFPOSX1 \Mem_reg[6][27]  ( .D(n2505), .CLK(clk), .Q(\Mem[6][27] ) );
  DFFPOSX1 \Mem_reg[6][26]  ( .D(n2504), .CLK(clk), .Q(\Mem[6][26] ) );
  DFFPOSX1 \Mem_reg[6][25]  ( .D(n2503), .CLK(clk), .Q(\Mem[6][25] ) );
  DFFPOSX1 \Mem_reg[6][24]  ( .D(n2502), .CLK(clk), .Q(\Mem[6][24] ) );
  DFFPOSX1 \Mem_reg[6][23]  ( .D(n2501), .CLK(clk), .Q(\Mem[6][23] ) );
  DFFPOSX1 \Mem_reg[6][22]  ( .D(n2500), .CLK(clk), .Q(\Mem[6][22] ) );
  DFFPOSX1 \Mem_reg[6][21]  ( .D(n2499), .CLK(clk), .Q(\Mem[6][21] ) );
  DFFPOSX1 \Mem_reg[6][20]  ( .D(n2498), .CLK(clk), .Q(\Mem[6][20] ) );
  DFFPOSX1 \Mem_reg[6][19]  ( .D(n2497), .CLK(clk), .Q(\Mem[6][19] ) );
  DFFPOSX1 \Mem_reg[6][18]  ( .D(n2496), .CLK(clk), .Q(\Mem[6][18] ) );
  DFFPOSX1 \Mem_reg[6][17]  ( .D(n2495), .CLK(clk), .Q(\Mem[6][17] ) );
  DFFPOSX1 \Mem_reg[6][16]  ( .D(n2494), .CLK(clk), .Q(\Mem[6][16] ) );
  DFFPOSX1 \Mem_reg[6][15]  ( .D(n2493), .CLK(clk), .Q(\Mem[6][15] ) );
  DFFPOSX1 \Mem_reg[6][14]  ( .D(n2492), .CLK(clk), .Q(\Mem[6][14] ) );
  DFFPOSX1 \Mem_reg[6][13]  ( .D(n2491), .CLK(clk), .Q(\Mem[6][13] ) );
  DFFPOSX1 \Mem_reg[6][12]  ( .D(n2490), .CLK(clk), .Q(\Mem[6][12] ) );
  DFFPOSX1 \Mem_reg[6][11]  ( .D(n2489), .CLK(clk), .Q(\Mem[6][11] ) );
  DFFPOSX1 \Mem_reg[6][10]  ( .D(n2488), .CLK(clk), .Q(\Mem[6][10] ) );
  DFFPOSX1 \Mem_reg[6][9]  ( .D(n2487), .CLK(clk), .Q(\Mem[6][9] ) );
  DFFPOSX1 \Mem_reg[6][8]  ( .D(n2486), .CLK(clk), .Q(\Mem[6][8] ) );
  DFFPOSX1 \Mem_reg[6][7]  ( .D(n2485), .CLK(clk), .Q(\Mem[6][7] ) );
  DFFPOSX1 \Mem_reg[6][6]  ( .D(n2484), .CLK(clk), .Q(\Mem[6][6] ) );
  DFFPOSX1 \Mem_reg[6][5]  ( .D(n2483), .CLK(clk), .Q(\Mem[6][5] ) );
  DFFPOSX1 \Mem_reg[6][4]  ( .D(n2482), .CLK(clk), .Q(\Mem[6][4] ) );
  DFFPOSX1 \Mem_reg[6][3]  ( .D(n2481), .CLK(clk), .Q(\Mem[6][3] ) );
  DFFPOSX1 \Mem_reg[6][2]  ( .D(n2480), .CLK(clk), .Q(\Mem[6][2] ) );
  DFFPOSX1 \Mem_reg[6][1]  ( .D(n2479), .CLK(clk), .Q(\Mem[6][1] ) );
  DFFPOSX1 \Mem_reg[6][0]  ( .D(n2478), .CLK(clk), .Q(\Mem[6][0] ) );
  DFFPOSX1 \Mem_reg[5][31]  ( .D(n2477), .CLK(clk), .Q(\Mem[5][31] ) );
  DFFPOSX1 \Mem_reg[5][30]  ( .D(n2476), .CLK(clk), .Q(\Mem[5][30] ) );
  DFFPOSX1 \Mem_reg[5][29]  ( .D(n2475), .CLK(clk), .Q(\Mem[5][29] ) );
  DFFPOSX1 \Mem_reg[5][28]  ( .D(n2474), .CLK(clk), .Q(\Mem[5][28] ) );
  DFFPOSX1 \Mem_reg[5][27]  ( .D(n2473), .CLK(clk), .Q(\Mem[5][27] ) );
  DFFPOSX1 \Mem_reg[5][26]  ( .D(n2472), .CLK(clk), .Q(\Mem[5][26] ) );
  DFFPOSX1 \Mem_reg[5][25]  ( .D(n2471), .CLK(clk), .Q(\Mem[5][25] ) );
  DFFPOSX1 \Mem_reg[5][24]  ( .D(n2470), .CLK(clk), .Q(\Mem[5][24] ) );
  DFFPOSX1 \Mem_reg[5][23]  ( .D(n2469), .CLK(clk), .Q(\Mem[5][23] ) );
  DFFPOSX1 \Mem_reg[5][22]  ( .D(n2468), .CLK(clk), .Q(\Mem[5][22] ) );
  DFFPOSX1 \Mem_reg[5][21]  ( .D(n2467), .CLK(clk), .Q(\Mem[5][21] ) );
  DFFPOSX1 \Mem_reg[5][20]  ( .D(n2466), .CLK(clk), .Q(\Mem[5][20] ) );
  DFFPOSX1 \Mem_reg[5][19]  ( .D(n2465), .CLK(clk), .Q(\Mem[5][19] ) );
  DFFPOSX1 \Mem_reg[5][18]  ( .D(n2464), .CLK(clk), .Q(\Mem[5][18] ) );
  DFFPOSX1 \Mem_reg[5][17]  ( .D(n2463), .CLK(clk), .Q(\Mem[5][17] ) );
  DFFPOSX1 \Mem_reg[5][16]  ( .D(n2462), .CLK(clk), .Q(\Mem[5][16] ) );
  DFFPOSX1 \Mem_reg[5][15]  ( .D(n2461), .CLK(clk), .Q(\Mem[5][15] ) );
  DFFPOSX1 \Mem_reg[5][14]  ( .D(n2460), .CLK(clk), .Q(\Mem[5][14] ) );
  DFFPOSX1 \Mem_reg[5][13]  ( .D(n2459), .CLK(clk), .Q(\Mem[5][13] ) );
  DFFPOSX1 \Mem_reg[5][12]  ( .D(n2458), .CLK(clk), .Q(\Mem[5][12] ) );
  DFFPOSX1 \Mem_reg[5][11]  ( .D(n2457), .CLK(clk), .Q(\Mem[5][11] ) );
  DFFPOSX1 \Mem_reg[5][10]  ( .D(n2456), .CLK(clk), .Q(\Mem[5][10] ) );
  DFFPOSX1 \Mem_reg[5][9]  ( .D(n2455), .CLK(clk), .Q(\Mem[5][9] ) );
  DFFPOSX1 \Mem_reg[5][8]  ( .D(n2454), .CLK(clk), .Q(\Mem[5][8] ) );
  DFFPOSX1 \Mem_reg[5][7]  ( .D(n2453), .CLK(clk), .Q(\Mem[5][7] ) );
  DFFPOSX1 \Mem_reg[5][6]  ( .D(n2452), .CLK(clk), .Q(\Mem[5][6] ) );
  DFFPOSX1 \Mem_reg[5][5]  ( .D(n2451), .CLK(clk), .Q(\Mem[5][5] ) );
  DFFPOSX1 \Mem_reg[5][4]  ( .D(n2450), .CLK(clk), .Q(\Mem[5][4] ) );
  DFFPOSX1 \Mem_reg[5][3]  ( .D(n2449), .CLK(clk), .Q(\Mem[5][3] ) );
  DFFPOSX1 \Mem_reg[5][2]  ( .D(n2448), .CLK(clk), .Q(\Mem[5][2] ) );
  DFFPOSX1 \Mem_reg[5][1]  ( .D(n2447), .CLK(clk), .Q(\Mem[5][1] ) );
  DFFPOSX1 \Mem_reg[5][0]  ( .D(n2446), .CLK(clk), .Q(\Mem[5][0] ) );
  DFFPOSX1 \Mem_reg[4][31]  ( .D(n2445), .CLK(clk), .Q(\Mem[4][31] ) );
  DFFPOSX1 \Mem_reg[4][30]  ( .D(n2444), .CLK(clk), .Q(\Mem[4][30] ) );
  DFFPOSX1 \Mem_reg[4][29]  ( .D(n2443), .CLK(clk), .Q(\Mem[4][29] ) );
  DFFPOSX1 \Mem_reg[4][28]  ( .D(n2442), .CLK(clk), .Q(\Mem[4][28] ) );
  DFFPOSX1 \Mem_reg[4][27]  ( .D(n2441), .CLK(clk), .Q(\Mem[4][27] ) );
  DFFPOSX1 \Mem_reg[4][26]  ( .D(n2440), .CLK(clk), .Q(\Mem[4][26] ) );
  DFFPOSX1 \Mem_reg[4][25]  ( .D(n2439), .CLK(clk), .Q(\Mem[4][25] ) );
  DFFPOSX1 \Mem_reg[4][24]  ( .D(n2438), .CLK(clk), .Q(\Mem[4][24] ) );
  DFFPOSX1 \Mem_reg[4][23]  ( .D(n2437), .CLK(clk), .Q(\Mem[4][23] ) );
  DFFPOSX1 \Mem_reg[4][22]  ( .D(n2436), .CLK(clk), .Q(\Mem[4][22] ) );
  DFFPOSX1 \Mem_reg[4][21]  ( .D(n2435), .CLK(clk), .Q(\Mem[4][21] ) );
  DFFPOSX1 \Mem_reg[4][20]  ( .D(n2434), .CLK(clk), .Q(\Mem[4][20] ) );
  DFFPOSX1 \Mem_reg[4][19]  ( .D(n2433), .CLK(clk), .Q(\Mem[4][19] ) );
  DFFPOSX1 \Mem_reg[4][18]  ( .D(n2432), .CLK(clk), .Q(\Mem[4][18] ) );
  DFFPOSX1 \Mem_reg[4][17]  ( .D(n2431), .CLK(clk), .Q(\Mem[4][17] ) );
  DFFPOSX1 \Mem_reg[4][16]  ( .D(n2430), .CLK(clk), .Q(\Mem[4][16] ) );
  DFFPOSX1 \Mem_reg[4][15]  ( .D(n2429), .CLK(clk), .Q(\Mem[4][15] ) );
  DFFPOSX1 \Mem_reg[4][14]  ( .D(n2428), .CLK(clk), .Q(\Mem[4][14] ) );
  DFFPOSX1 \Mem_reg[4][13]  ( .D(n2427), .CLK(clk), .Q(\Mem[4][13] ) );
  DFFPOSX1 \Mem_reg[4][12]  ( .D(n2426), .CLK(clk), .Q(\Mem[4][12] ) );
  DFFPOSX1 \Mem_reg[4][11]  ( .D(n2425), .CLK(clk), .Q(\Mem[4][11] ) );
  DFFPOSX1 \Mem_reg[4][10]  ( .D(n2424), .CLK(clk), .Q(\Mem[4][10] ) );
  DFFPOSX1 \Mem_reg[4][9]  ( .D(n2423), .CLK(clk), .Q(\Mem[4][9] ) );
  DFFPOSX1 \Mem_reg[4][8]  ( .D(n2422), .CLK(clk), .Q(\Mem[4][8] ) );
  DFFPOSX1 \Mem_reg[4][7]  ( .D(n2421), .CLK(clk), .Q(\Mem[4][7] ) );
  DFFPOSX1 \Mem_reg[4][6]  ( .D(n2420), .CLK(clk), .Q(\Mem[4][6] ) );
  DFFPOSX1 \Mem_reg[4][5]  ( .D(n2419), .CLK(clk), .Q(\Mem[4][5] ) );
  DFFPOSX1 \Mem_reg[4][4]  ( .D(n2418), .CLK(clk), .Q(\Mem[4][4] ) );
  DFFPOSX1 \Mem_reg[4][3]  ( .D(n2417), .CLK(clk), .Q(\Mem[4][3] ) );
  DFFPOSX1 \Mem_reg[4][2]  ( .D(n2416), .CLK(clk), .Q(\Mem[4][2] ) );
  DFFPOSX1 \Mem_reg[4][1]  ( .D(n2415), .CLK(clk), .Q(\Mem[4][1] ) );
  DFFPOSX1 \Mem_reg[4][0]  ( .D(n2414), .CLK(clk), .Q(\Mem[4][0] ) );
  DFFPOSX1 \Mem_reg[3][31]  ( .D(n2413), .CLK(clk), .Q(\Mem[3][31] ) );
  DFFPOSX1 \Mem_reg[3][30]  ( .D(n2412), .CLK(clk), .Q(\Mem[3][30] ) );
  DFFPOSX1 \Mem_reg[3][29]  ( .D(n2411), .CLK(clk), .Q(\Mem[3][29] ) );
  DFFPOSX1 \Mem_reg[3][28]  ( .D(n2410), .CLK(clk), .Q(\Mem[3][28] ) );
  DFFPOSX1 \Mem_reg[3][27]  ( .D(n2409), .CLK(clk), .Q(\Mem[3][27] ) );
  DFFPOSX1 \Mem_reg[3][26]  ( .D(n2408), .CLK(clk), .Q(\Mem[3][26] ) );
  DFFPOSX1 \Mem_reg[3][25]  ( .D(n2407), .CLK(clk), .Q(\Mem[3][25] ) );
  DFFPOSX1 \Mem_reg[3][24]  ( .D(n2406), .CLK(clk), .Q(\Mem[3][24] ) );
  DFFPOSX1 \Mem_reg[3][23]  ( .D(n2405), .CLK(clk), .Q(\Mem[3][23] ) );
  DFFPOSX1 \Mem_reg[3][22]  ( .D(n2404), .CLK(clk), .Q(\Mem[3][22] ) );
  DFFPOSX1 \Mem_reg[3][21]  ( .D(n2403), .CLK(clk), .Q(\Mem[3][21] ) );
  DFFPOSX1 \Mem_reg[3][20]  ( .D(n2402), .CLK(clk), .Q(\Mem[3][20] ) );
  DFFPOSX1 \Mem_reg[3][19]  ( .D(n2401), .CLK(clk), .Q(\Mem[3][19] ) );
  DFFPOSX1 \Mem_reg[3][18]  ( .D(n2400), .CLK(clk), .Q(\Mem[3][18] ) );
  DFFPOSX1 \Mem_reg[3][17]  ( .D(n2399), .CLK(clk), .Q(\Mem[3][17] ) );
  DFFPOSX1 \Mem_reg[3][16]  ( .D(n2398), .CLK(clk), .Q(\Mem[3][16] ) );
  DFFPOSX1 \Mem_reg[3][15]  ( .D(n2397), .CLK(clk), .Q(\Mem[3][15] ) );
  DFFPOSX1 \Mem_reg[3][14]  ( .D(n2396), .CLK(clk), .Q(\Mem[3][14] ) );
  DFFPOSX1 \Mem_reg[3][13]  ( .D(n2395), .CLK(clk), .Q(\Mem[3][13] ) );
  DFFPOSX1 \Mem_reg[3][12]  ( .D(n2394), .CLK(clk), .Q(\Mem[3][12] ) );
  DFFPOSX1 \Mem_reg[3][11]  ( .D(n2393), .CLK(clk), .Q(\Mem[3][11] ) );
  DFFPOSX1 \Mem_reg[3][10]  ( .D(n2392), .CLK(clk), .Q(\Mem[3][10] ) );
  DFFPOSX1 \Mem_reg[3][9]  ( .D(n2391), .CLK(clk), .Q(\Mem[3][9] ) );
  DFFPOSX1 \Mem_reg[3][8]  ( .D(n2390), .CLK(clk), .Q(\Mem[3][8] ) );
  DFFPOSX1 \Mem_reg[3][7]  ( .D(n2389), .CLK(clk), .Q(\Mem[3][7] ) );
  DFFPOSX1 \Mem_reg[3][6]  ( .D(n2388), .CLK(clk), .Q(\Mem[3][6] ) );
  DFFPOSX1 \Mem_reg[3][5]  ( .D(n2387), .CLK(clk), .Q(\Mem[3][5] ) );
  DFFPOSX1 \Mem_reg[3][4]  ( .D(n2386), .CLK(clk), .Q(\Mem[3][4] ) );
  DFFPOSX1 \Mem_reg[3][3]  ( .D(n2385), .CLK(clk), .Q(\Mem[3][3] ) );
  DFFPOSX1 \Mem_reg[3][2]  ( .D(n2384), .CLK(clk), .Q(\Mem[3][2] ) );
  DFFPOSX1 \Mem_reg[3][1]  ( .D(n2383), .CLK(clk), .Q(\Mem[3][1] ) );
  DFFPOSX1 \Mem_reg[3][0]  ( .D(n2382), .CLK(clk), .Q(\Mem[3][0] ) );
  DFFPOSX1 \Mem_reg[2][31]  ( .D(n2381), .CLK(clk), .Q(\Mem[2][31] ) );
  DFFPOSX1 \Mem_reg[2][30]  ( .D(n2380), .CLK(clk), .Q(\Mem[2][30] ) );
  DFFPOSX1 \Mem_reg[2][29]  ( .D(n2379), .CLK(clk), .Q(\Mem[2][29] ) );
  DFFPOSX1 \Mem_reg[2][28]  ( .D(n2378), .CLK(clk), .Q(\Mem[2][28] ) );
  DFFPOSX1 \Mem_reg[2][27]  ( .D(n2377), .CLK(clk), .Q(\Mem[2][27] ) );
  DFFPOSX1 \Mem_reg[2][26]  ( .D(n2376), .CLK(clk), .Q(\Mem[2][26] ) );
  DFFPOSX1 \Mem_reg[2][25]  ( .D(n2375), .CLK(clk), .Q(\Mem[2][25] ) );
  DFFPOSX1 \Mem_reg[2][24]  ( .D(n2374), .CLK(clk), .Q(\Mem[2][24] ) );
  DFFPOSX1 \Mem_reg[2][23]  ( .D(n2373), .CLK(clk), .Q(\Mem[2][23] ) );
  DFFPOSX1 \Mem_reg[2][22]  ( .D(n2372), .CLK(clk), .Q(\Mem[2][22] ) );
  DFFPOSX1 \Mem_reg[2][21]  ( .D(n2371), .CLK(clk), .Q(\Mem[2][21] ) );
  DFFPOSX1 \Mem_reg[2][20]  ( .D(n2370), .CLK(clk), .Q(\Mem[2][20] ) );
  DFFPOSX1 \Mem_reg[2][19]  ( .D(n2369), .CLK(clk), .Q(\Mem[2][19] ) );
  DFFPOSX1 \Mem_reg[2][18]  ( .D(n2368), .CLK(clk), .Q(\Mem[2][18] ) );
  DFFPOSX1 \Mem_reg[2][17]  ( .D(n2367), .CLK(clk), .Q(\Mem[2][17] ) );
  DFFPOSX1 \Mem_reg[2][16]  ( .D(n2366), .CLK(clk), .Q(\Mem[2][16] ) );
  DFFPOSX1 \Mem_reg[2][15]  ( .D(n2365), .CLK(clk), .Q(\Mem[2][15] ) );
  DFFPOSX1 \Mem_reg[2][14]  ( .D(n2364), .CLK(clk), .Q(\Mem[2][14] ) );
  DFFPOSX1 \Mem_reg[2][13]  ( .D(n2363), .CLK(clk), .Q(\Mem[2][13] ) );
  DFFPOSX1 \Mem_reg[2][12]  ( .D(n2362), .CLK(clk), .Q(\Mem[2][12] ) );
  DFFPOSX1 \Mem_reg[2][11]  ( .D(n2361), .CLK(clk), .Q(\Mem[2][11] ) );
  DFFPOSX1 \Mem_reg[2][10]  ( .D(n2360), .CLK(clk), .Q(\Mem[2][10] ) );
  DFFPOSX1 \Mem_reg[2][9]  ( .D(n2359), .CLK(clk), .Q(\Mem[2][9] ) );
  DFFPOSX1 \Mem_reg[2][8]  ( .D(n2358), .CLK(clk), .Q(\Mem[2][8] ) );
  DFFPOSX1 \Mem_reg[2][7]  ( .D(n2357), .CLK(clk), .Q(\Mem[2][7] ) );
  DFFPOSX1 \Mem_reg[2][6]  ( .D(n2356), .CLK(clk), .Q(\Mem[2][6] ) );
  DFFPOSX1 \Mem_reg[2][5]  ( .D(n2355), .CLK(clk), .Q(\Mem[2][5] ) );
  DFFPOSX1 \Mem_reg[2][4]  ( .D(n2354), .CLK(clk), .Q(\Mem[2][4] ) );
  DFFPOSX1 \Mem_reg[2][3]  ( .D(n2353), .CLK(clk), .Q(\Mem[2][3] ) );
  DFFPOSX1 \Mem_reg[2][2]  ( .D(n2352), .CLK(clk), .Q(\Mem[2][2] ) );
  DFFPOSX1 \Mem_reg[2][1]  ( .D(n2351), .CLK(clk), .Q(\Mem[2][1] ) );
  DFFPOSX1 \Mem_reg[2][0]  ( .D(n2350), .CLK(clk), .Q(\Mem[2][0] ) );
  DFFPOSX1 \Mem_reg[1][31]  ( .D(n2349), .CLK(clk), .Q(\Mem[1][31] ) );
  DFFPOSX1 \Mem_reg[1][30]  ( .D(n2348), .CLK(clk), .Q(\Mem[1][30] ) );
  DFFPOSX1 \Mem_reg[1][29]  ( .D(n2347), .CLK(clk), .Q(\Mem[1][29] ) );
  DFFPOSX1 \Mem_reg[1][28]  ( .D(n2346), .CLK(clk), .Q(\Mem[1][28] ) );
  DFFPOSX1 \Mem_reg[1][27]  ( .D(n2345), .CLK(clk), .Q(\Mem[1][27] ) );
  DFFPOSX1 \Mem_reg[1][26]  ( .D(n2344), .CLK(clk), .Q(\Mem[1][26] ) );
  DFFPOSX1 \Mem_reg[1][25]  ( .D(n2343), .CLK(clk), .Q(\Mem[1][25] ) );
  DFFPOSX1 \Mem_reg[1][24]  ( .D(n2342), .CLK(clk), .Q(\Mem[1][24] ) );
  DFFPOSX1 \Mem_reg[1][23]  ( .D(n2341), .CLK(clk), .Q(\Mem[1][23] ) );
  DFFPOSX1 \Mem_reg[1][22]  ( .D(n2340), .CLK(clk), .Q(\Mem[1][22] ) );
  DFFPOSX1 \Mem_reg[1][21]  ( .D(n2339), .CLK(clk), .Q(\Mem[1][21] ) );
  DFFPOSX1 \Mem_reg[1][20]  ( .D(n2338), .CLK(clk), .Q(\Mem[1][20] ) );
  DFFPOSX1 \Mem_reg[1][19]  ( .D(n2337), .CLK(clk), .Q(\Mem[1][19] ) );
  DFFPOSX1 \Mem_reg[1][18]  ( .D(n2336), .CLK(clk), .Q(\Mem[1][18] ) );
  DFFPOSX1 \Mem_reg[1][17]  ( .D(n2335), .CLK(clk), .Q(\Mem[1][17] ) );
  DFFPOSX1 \Mem_reg[1][16]  ( .D(n2334), .CLK(clk), .Q(\Mem[1][16] ) );
  DFFPOSX1 \Mem_reg[1][15]  ( .D(n2333), .CLK(clk), .Q(\Mem[1][15] ) );
  DFFPOSX1 \Mem_reg[1][14]  ( .D(n2332), .CLK(clk), .Q(\Mem[1][14] ) );
  DFFPOSX1 \Mem_reg[1][13]  ( .D(n2331), .CLK(clk), .Q(\Mem[1][13] ) );
  DFFPOSX1 \Mem_reg[1][12]  ( .D(n2330), .CLK(clk), .Q(\Mem[1][12] ) );
  DFFPOSX1 \Mem_reg[1][11]  ( .D(n2329), .CLK(clk), .Q(\Mem[1][11] ) );
  DFFPOSX1 \Mem_reg[1][10]  ( .D(n2328), .CLK(clk), .Q(\Mem[1][10] ) );
  DFFPOSX1 \Mem_reg[1][9]  ( .D(n2327), .CLK(clk), .Q(\Mem[1][9] ) );
  DFFPOSX1 \Mem_reg[1][8]  ( .D(n2326), .CLK(clk), .Q(\Mem[1][8] ) );
  DFFPOSX1 \Mem_reg[1][7]  ( .D(n2325), .CLK(clk), .Q(\Mem[1][7] ) );
  DFFPOSX1 \Mem_reg[1][6]  ( .D(n2324), .CLK(clk), .Q(\Mem[1][6] ) );
  DFFPOSX1 \Mem_reg[1][5]  ( .D(n2323), .CLK(clk), .Q(\Mem[1][5] ) );
  DFFPOSX1 \Mem_reg[1][4]  ( .D(n2322), .CLK(clk), .Q(\Mem[1][4] ) );
  DFFPOSX1 \Mem_reg[1][3]  ( .D(n2321), .CLK(clk), .Q(\Mem[1][3] ) );
  DFFPOSX1 \Mem_reg[1][2]  ( .D(n2320), .CLK(clk), .Q(\Mem[1][2] ) );
  DFFPOSX1 \Mem_reg[1][1]  ( .D(n2319), .CLK(clk), .Q(\Mem[1][1] ) );
  DFFPOSX1 \Mem_reg[1][0]  ( .D(n2318), .CLK(clk), .Q(\Mem[1][0] ) );
  DFFPOSX1 \Mem_reg[0][31]  ( .D(n2317), .CLK(clk), .Q(\Mem[0][31] ) );
  DFFPOSX1 \Mem_reg[0][30]  ( .D(n2316), .CLK(clk), .Q(\Mem[0][30] ) );
  DFFPOSX1 \Mem_reg[0][29]  ( .D(n2315), .CLK(clk), .Q(\Mem[0][29] ) );
  DFFPOSX1 \Mem_reg[0][28]  ( .D(n2314), .CLK(clk), .Q(\Mem[0][28] ) );
  DFFPOSX1 \Mem_reg[0][27]  ( .D(n2313), .CLK(clk), .Q(\Mem[0][27] ) );
  DFFPOSX1 \Mem_reg[0][26]  ( .D(n2312), .CLK(clk), .Q(\Mem[0][26] ) );
  DFFPOSX1 \Mem_reg[0][25]  ( .D(n2311), .CLK(clk), .Q(\Mem[0][25] ) );
  DFFPOSX1 \Mem_reg[0][24]  ( .D(n2310), .CLK(clk), .Q(\Mem[0][24] ) );
  DFFPOSX1 \Mem_reg[0][23]  ( .D(n2309), .CLK(clk), .Q(\Mem[0][23] ) );
  DFFPOSX1 \Mem_reg[0][22]  ( .D(n2308), .CLK(clk), .Q(\Mem[0][22] ) );
  DFFPOSX1 \Mem_reg[0][21]  ( .D(n2307), .CLK(clk), .Q(\Mem[0][21] ) );
  DFFPOSX1 \Mem_reg[0][20]  ( .D(n2306), .CLK(clk), .Q(\Mem[0][20] ) );
  DFFPOSX1 \Mem_reg[0][19]  ( .D(n2305), .CLK(clk), .Q(\Mem[0][19] ) );
  DFFPOSX1 \Mem_reg[0][18]  ( .D(n2304), .CLK(clk), .Q(\Mem[0][18] ) );
  DFFPOSX1 \Mem_reg[0][17]  ( .D(n2303), .CLK(clk), .Q(\Mem[0][17] ) );
  DFFPOSX1 \Mem_reg[0][16]  ( .D(n2302), .CLK(clk), .Q(\Mem[0][16] ) );
  DFFPOSX1 \Mem_reg[0][15]  ( .D(n2301), .CLK(clk), .Q(\Mem[0][15] ) );
  DFFPOSX1 \Mem_reg[0][14]  ( .D(n2300), .CLK(clk), .Q(\Mem[0][14] ) );
  DFFPOSX1 \Mem_reg[0][13]  ( .D(n2299), .CLK(clk), .Q(\Mem[0][13] ) );
  DFFPOSX1 \Mem_reg[0][12]  ( .D(n2298), .CLK(clk), .Q(\Mem[0][12] ) );
  DFFPOSX1 \Mem_reg[0][11]  ( .D(n2297), .CLK(clk), .Q(\Mem[0][11] ) );
  DFFPOSX1 \Mem_reg[0][10]  ( .D(n2296), .CLK(clk), .Q(\Mem[0][10] ) );
  DFFPOSX1 \Mem_reg[0][9]  ( .D(n2295), .CLK(clk), .Q(\Mem[0][9] ) );
  DFFPOSX1 \Mem_reg[0][8]  ( .D(n2294), .CLK(clk), .Q(\Mem[0][8] ) );
  DFFPOSX1 \Mem_reg[0][7]  ( .D(n2293), .CLK(clk), .Q(\Mem[0][7] ) );
  DFFPOSX1 \Mem_reg[0][6]  ( .D(n2292), .CLK(clk), .Q(\Mem[0][6] ) );
  DFFPOSX1 \Mem_reg[0][5]  ( .D(n2291), .CLK(clk), .Q(\Mem[0][5] ) );
  DFFPOSX1 \Mem_reg[0][4]  ( .D(n2290), .CLK(clk), .Q(\Mem[0][4] ) );
  DFFPOSX1 \Mem_reg[0][3]  ( .D(n2289), .CLK(clk), .Q(\Mem[0][3] ) );
  DFFPOSX1 \Mem_reg[0][2]  ( .D(n2288), .CLK(clk), .Q(\Mem[0][2] ) );
  DFFPOSX1 \Mem_reg[0][1]  ( .D(n2287), .CLK(clk), .Q(\Mem[0][1] ) );
  DFFPOSX1 \Mem_reg[0][0]  ( .D(n2286), .CLK(clk), .Q(\Mem[0][0] ) );
  OAI21X1 U2 ( .A(n6925), .B(n6554), .C(n3), .Y(n2497) );
  NAND2X1 U3 ( .A(\Mem[6][19] ), .B(n6928), .Y(n3) );
  OAI21X1 U4 ( .A(n6924), .B(n6544), .C(n5), .Y(n2498) );
  NAND2X1 U5 ( .A(\Mem[6][20] ), .B(n6928), .Y(n5) );
  OAI21X1 U6 ( .A(n6924), .B(n6539), .C(n7), .Y(n2499) );
  NAND2X1 U7 ( .A(\Mem[6][21] ), .B(n6928), .Y(n7) );
  OAI21X1 U8 ( .A(n6924), .B(n6534), .C(n9), .Y(n2500) );
  NAND2X1 U9 ( .A(\Mem[6][22] ), .B(n6927), .Y(n9) );
  OAI21X1 U10 ( .A(n6924), .B(n6529), .C(n11), .Y(n2501) );
  NAND2X1 U11 ( .A(\Mem[6][23] ), .B(n6927), .Y(n11) );
  OAI21X1 U12 ( .A(n6924), .B(n6524), .C(n13), .Y(n2502) );
  NAND2X1 U13 ( .A(\Mem[6][24] ), .B(n6927), .Y(n13) );
  OAI21X1 U14 ( .A(n6924), .B(n6519), .C(n15), .Y(n2503) );
  NAND2X1 U15 ( .A(\Mem[6][25] ), .B(n6927), .Y(n15) );
  OAI21X1 U16 ( .A(n6924), .B(n6514), .C(n17), .Y(n2504) );
  NAND2X1 U17 ( .A(\Mem[6][26] ), .B(n6927), .Y(n17) );
  OAI21X1 U18 ( .A(n6924), .B(n6509), .C(n19), .Y(n2505) );
  NAND2X1 U19 ( .A(\Mem[6][27] ), .B(n6927), .Y(n19) );
  OAI21X1 U20 ( .A(n6924), .B(n6504), .C(n21), .Y(n2506) );
  NAND2X1 U21 ( .A(\Mem[6][28] ), .B(n6927), .Y(n21) );
  OAI21X1 U22 ( .A(n6924), .B(n6499), .C(n23), .Y(n2507) );
  NAND2X1 U23 ( .A(\Mem[6][29] ), .B(n6927), .Y(n23) );
  OAI21X1 U24 ( .A(n6924), .B(n6489), .C(n25), .Y(n2508) );
  NAND2X1 U25 ( .A(\Mem[6][30] ), .B(n6927), .Y(n25) );
  OAI21X1 U26 ( .A(n6924), .B(n6484), .C(n27), .Y(n2509) );
  NAND2X1 U27 ( .A(\Mem[6][31] ), .B(n6927), .Y(n27) );
  OAI21X1 U28 ( .A(n6921), .B(n6604), .C(n30), .Y(n2510) );
  NAND2X1 U29 ( .A(\Mem[7][0] ), .B(n6923), .Y(n30) );
  OAI21X1 U30 ( .A(n6920), .B(n6549), .C(n32), .Y(n2511) );
  NAND2X1 U31 ( .A(\Mem[7][1] ), .B(n6923), .Y(n32) );
  OAI21X1 U32 ( .A(n6920), .B(n6494), .C(n34), .Y(n2512) );
  NAND2X1 U33 ( .A(\Mem[7][2] ), .B(n6922), .Y(n34) );
  OAI21X1 U34 ( .A(n6920), .B(n6479), .C(n36), .Y(n2513) );
  NAND2X1 U35 ( .A(\Mem[7][3] ), .B(n6922), .Y(n36) );
  OAI21X1 U36 ( .A(n6920), .B(n6474), .C(n38), .Y(n2514) );
  NAND2X1 U37 ( .A(\Mem[7][4] ), .B(n6922), .Y(n38) );
  OAI21X1 U38 ( .A(n6920), .B(n6469), .C(n40), .Y(n2515) );
  NAND2X1 U39 ( .A(\Mem[7][5] ), .B(n6922), .Y(n40) );
  OAI21X1 U40 ( .A(n6920), .B(n6464), .C(n42), .Y(n2516) );
  NAND2X1 U41 ( .A(\Mem[7][6] ), .B(n6922), .Y(n42) );
  OAI21X1 U42 ( .A(n6920), .B(n6459), .C(n44), .Y(n2517) );
  NAND2X1 U43 ( .A(\Mem[7][7] ), .B(n6922), .Y(n44) );
  OAI21X1 U44 ( .A(n6920), .B(n6454), .C(n46), .Y(n2518) );
  NAND2X1 U45 ( .A(\Mem[7][8] ), .B(n6922), .Y(n46) );
  OAI21X1 U46 ( .A(n6920), .B(n6449), .C(n48), .Y(n2519) );
  NAND2X1 U47 ( .A(\Mem[7][9] ), .B(n6922), .Y(n48) );
  OAI21X1 U48 ( .A(n6920), .B(n6599), .C(n50), .Y(n2520) );
  NAND2X1 U49 ( .A(\Mem[7][10] ), .B(n6922), .Y(n50) );
  OAI21X1 U50 ( .A(n6920), .B(n6594), .C(n52), .Y(n2521) );
  NAND2X1 U51 ( .A(\Mem[7][11] ), .B(n6922), .Y(n52) );
  OAI21X1 U52 ( .A(n6920), .B(n6589), .C(n54), .Y(n2522) );
  NAND2X1 U53 ( .A(\Mem[7][12] ), .B(n6921), .Y(n54) );
  OAI21X1 U54 ( .A(n6921), .B(n6584), .C(n56), .Y(n2523) );
  NAND2X1 U55 ( .A(\Mem[7][13] ), .B(n6921), .Y(n56) );
  OAI21X1 U56 ( .A(n6921), .B(n6579), .C(n58), .Y(n2524) );
  NAND2X1 U57 ( .A(\Mem[7][14] ), .B(n6921), .Y(n58) );
  OAI21X1 U58 ( .A(n6921), .B(n6574), .C(n60), .Y(n2525) );
  NAND2X1 U59 ( .A(\Mem[7][15] ), .B(n6921), .Y(n60) );
  OAI21X1 U60 ( .A(n6921), .B(n6569), .C(n62), .Y(n2526) );
  NAND2X1 U61 ( .A(\Mem[7][16] ), .B(n6921), .Y(n62) );
  OAI21X1 U62 ( .A(n6921), .B(n6564), .C(n64), .Y(n2527) );
  NAND2X1 U63 ( .A(\Mem[7][17] ), .B(n6921), .Y(n64) );
  OAI21X1 U64 ( .A(n6921), .B(n6559), .C(n66), .Y(n2528) );
  NAND2X1 U65 ( .A(\Mem[7][18] ), .B(n6921), .Y(n66) );
  OAI21X1 U66 ( .A(n6554), .B(n6920), .C(n67), .Y(n2529) );
  NAND2X1 U67 ( .A(\Mem[7][19] ), .B(n6921), .Y(n67) );
  OAI21X1 U68 ( .A(n6544), .B(n6919), .C(n68), .Y(n2530) );
  NAND2X1 U69 ( .A(\Mem[7][20] ), .B(n6922), .Y(n68) );
  OAI21X1 U70 ( .A(n6539), .B(n6919), .C(n69), .Y(n2531) );
  NAND2X1 U71 ( .A(\Mem[7][21] ), .B(n6922), .Y(n69) );
  OAI21X1 U72 ( .A(n6534), .B(n6919), .C(n70), .Y(n2532) );
  NAND2X1 U73 ( .A(\Mem[7][22] ), .B(n6922), .Y(n70) );
  OAI21X1 U74 ( .A(n6529), .B(n6919), .C(n71), .Y(n2533) );
  NAND2X1 U75 ( .A(\Mem[7][23] ), .B(n6922), .Y(n71) );
  OAI21X1 U76 ( .A(n6524), .B(n6919), .C(n72), .Y(n2534) );
  NAND2X1 U77 ( .A(\Mem[7][24] ), .B(n6922), .Y(n72) );
  OAI21X1 U78 ( .A(n6519), .B(n6919), .C(n73), .Y(n2535) );
  NAND2X1 U79 ( .A(\Mem[7][25] ), .B(n6922), .Y(n73) );
  OAI21X1 U80 ( .A(n6514), .B(n6919), .C(n74), .Y(n2536) );
  NAND2X1 U81 ( .A(\Mem[7][26] ), .B(n6922), .Y(n74) );
  OAI21X1 U82 ( .A(n6509), .B(n6919), .C(n75), .Y(n2537) );
  NAND2X1 U83 ( .A(\Mem[7][27] ), .B(n6922), .Y(n75) );
  OAI21X1 U84 ( .A(n6504), .B(n6919), .C(n76), .Y(n2538) );
  NAND2X1 U85 ( .A(\Mem[7][28] ), .B(n6922), .Y(n76) );
  OAI21X1 U86 ( .A(n6499), .B(n6919), .C(n77), .Y(n2539) );
  NAND2X1 U87 ( .A(\Mem[7][29] ), .B(n6923), .Y(n77) );
  OAI21X1 U88 ( .A(n6489), .B(n6919), .C(n78), .Y(n2540) );
  NAND2X1 U89 ( .A(\Mem[7][30] ), .B(n6923), .Y(n78) );
  OAI21X1 U90 ( .A(n6484), .B(n6919), .C(n79), .Y(n2541) );
  NAND2X1 U91 ( .A(\Mem[7][31] ), .B(n6923), .Y(n79) );
  NAND2X1 U92 ( .A(n7021), .B(n7004), .Y(n28) );
  OAI21X1 U93 ( .A(n6604), .B(n6915), .C(n83), .Y(n2542) );
  NAND2X1 U94 ( .A(\Mem[8][0] ), .B(n6918), .Y(n83) );
  OAI21X1 U95 ( .A(n6549), .B(n6914), .C(n84), .Y(n2543) );
  NAND2X1 U96 ( .A(\Mem[8][1] ), .B(n6918), .Y(n84) );
  OAI21X1 U97 ( .A(n6494), .B(n6914), .C(n85), .Y(n2544) );
  NAND2X1 U98 ( .A(\Mem[8][2] ), .B(n6918), .Y(n85) );
  OAI21X1 U99 ( .A(n6479), .B(n6914), .C(n86), .Y(n2545) );
  NAND2X1 U100 ( .A(\Mem[8][3] ), .B(n6917), .Y(n86) );
  OAI21X1 U101 ( .A(n6474), .B(n6914), .C(n87), .Y(n2546) );
  NAND2X1 U102 ( .A(\Mem[8][4] ), .B(n6918), .Y(n87) );
  OAI21X1 U103 ( .A(n6469), .B(n6914), .C(n88), .Y(n2547) );
  NAND2X1 U104 ( .A(\Mem[8][5] ), .B(n6917), .Y(n88) );
  OAI21X1 U105 ( .A(n6464), .B(n6914), .C(n89), .Y(n2548) );
  NAND2X1 U106 ( .A(\Mem[8][6] ), .B(n6917), .Y(n89) );
  OAI21X1 U107 ( .A(n6459), .B(n6914), .C(n90), .Y(n2549) );
  NAND2X1 U108 ( .A(\Mem[8][7] ), .B(n6917), .Y(n90) );
  OAI21X1 U109 ( .A(n6454), .B(n6914), .C(n91), .Y(n2550) );
  NAND2X1 U110 ( .A(\Mem[8][8] ), .B(n6917), .Y(n91) );
  OAI21X1 U111 ( .A(n6449), .B(n6914), .C(n92), .Y(n2551) );
  NAND2X1 U112 ( .A(\Mem[8][9] ), .B(n6917), .Y(n92) );
  OAI21X1 U113 ( .A(n6599), .B(n6914), .C(n93), .Y(n2552) );
  NAND2X1 U114 ( .A(\Mem[8][10] ), .B(n6917), .Y(n93) );
  OAI21X1 U115 ( .A(n6594), .B(n6914), .C(n94), .Y(n2553) );
  NAND2X1 U116 ( .A(\Mem[8][11] ), .B(n6917), .Y(n94) );
  OAI21X1 U117 ( .A(n6589), .B(n6914), .C(n95), .Y(n2554) );
  NAND2X1 U118 ( .A(\Mem[8][12] ), .B(n6917), .Y(n95) );
  OAI21X1 U119 ( .A(n6584), .B(n6915), .C(n96), .Y(n2555) );
  NAND2X1 U120 ( .A(\Mem[8][13] ), .B(n6917), .Y(n96) );
  OAI21X1 U121 ( .A(n6579), .B(n6915), .C(n97), .Y(n2556) );
  NAND2X1 U122 ( .A(\Mem[8][14] ), .B(n6917), .Y(n97) );
  OAI21X1 U123 ( .A(n6574), .B(n6915), .C(n98), .Y(n2557) );
  NAND2X1 U124 ( .A(\Mem[8][15] ), .B(n6916), .Y(n98) );
  OAI21X1 U125 ( .A(n6569), .B(n6915), .C(n99), .Y(n2558) );
  NAND2X1 U126 ( .A(\Mem[8][16] ), .B(n6917), .Y(n99) );
  OAI21X1 U127 ( .A(n6564), .B(n6915), .C(n100), .Y(n2559) );
  NAND2X1 U128 ( .A(\Mem[8][17] ), .B(n6916), .Y(n100) );
  OAI21X1 U129 ( .A(n6559), .B(n6915), .C(n101), .Y(n2560) );
  NAND2X1 U130 ( .A(\Mem[8][18] ), .B(n6916), .Y(n101) );
  OAI21X1 U131 ( .A(n6554), .B(n6915), .C(n102), .Y(n2561) );
  NAND2X1 U132 ( .A(\Mem[8][19] ), .B(n6916), .Y(n102) );
  OAI21X1 U133 ( .A(n6544), .B(n6915), .C(n103), .Y(n2562) );
  NAND2X1 U134 ( .A(\Mem[8][20] ), .B(n6916), .Y(n103) );
  OAI21X1 U135 ( .A(n6539), .B(n6915), .C(n104), .Y(n2563) );
  NAND2X1 U136 ( .A(\Mem[8][21] ), .B(n6916), .Y(n104) );
  OAI21X1 U137 ( .A(n6534), .B(n6915), .C(n105), .Y(n2564) );
  NAND2X1 U138 ( .A(\Mem[8][22] ), .B(n6917), .Y(n105) );
  OAI21X1 U139 ( .A(n6529), .B(n6916), .C(n106), .Y(n2565) );
  NAND2X1 U140 ( .A(\Mem[8][23] ), .B(n6916), .Y(n106) );
  OAI21X1 U141 ( .A(n6524), .B(n6915), .C(n107), .Y(n2566) );
  NAND2X1 U142 ( .A(\Mem[8][24] ), .B(n6917), .Y(n107) );
  OAI21X1 U143 ( .A(n6519), .B(n6916), .C(n108), .Y(n2567) );
  NAND2X1 U144 ( .A(\Mem[8][25] ), .B(n6917), .Y(n108) );
  OAI21X1 U145 ( .A(n6514), .B(n6916), .C(n109), .Y(n2568) );
  NAND2X1 U146 ( .A(\Mem[8][26] ), .B(n6917), .Y(n109) );
  OAI21X1 U147 ( .A(n6509), .B(n6916), .C(n110), .Y(n2569) );
  NAND2X1 U148 ( .A(\Mem[8][27] ), .B(n6917), .Y(n110) );
  OAI21X1 U149 ( .A(n6504), .B(n6916), .C(n111), .Y(n2570) );
  NAND2X1 U150 ( .A(\Mem[8][28] ), .B(n6917), .Y(n111) );
  OAI21X1 U151 ( .A(n6499), .B(n6916), .C(n112), .Y(n2571) );
  NAND2X1 U152 ( .A(\Mem[8][29] ), .B(n6917), .Y(n112) );
  OAI21X1 U153 ( .A(n6489), .B(n6916), .C(n113), .Y(n2572) );
  NAND2X1 U154 ( .A(\Mem[8][30] ), .B(n6918), .Y(n113) );
  OAI21X1 U155 ( .A(n6484), .B(n6916), .C(n114), .Y(n2573) );
  NAND2X1 U156 ( .A(\Mem[8][31] ), .B(n6918), .Y(n114) );
  NAND2X1 U157 ( .A(n7016), .B(n7007), .Y(n82) );
  OAI21X1 U158 ( .A(n6605), .B(n6910), .C(n118), .Y(n2574) );
  NAND2X1 U159 ( .A(\Mem[9][0] ), .B(n6913), .Y(n118) );
  OAI21X1 U160 ( .A(n6550), .B(n6909), .C(n119), .Y(n2575) );
  NAND2X1 U161 ( .A(\Mem[9][1] ), .B(n6913), .Y(n119) );
  OAI21X1 U162 ( .A(n6495), .B(n6909), .C(n120), .Y(n2576) );
  NAND2X1 U163 ( .A(\Mem[9][2] ), .B(n6913), .Y(n120) );
  OAI21X1 U164 ( .A(n6480), .B(n6909), .C(n121), .Y(n2577) );
  NAND2X1 U165 ( .A(\Mem[9][3] ), .B(n6912), .Y(n121) );
  OAI21X1 U166 ( .A(n6475), .B(n6909), .C(n122), .Y(n2578) );
  NAND2X1 U167 ( .A(\Mem[9][4] ), .B(n6913), .Y(n122) );
  OAI21X1 U168 ( .A(n6470), .B(n6909), .C(n123), .Y(n2579) );
  NAND2X1 U169 ( .A(\Mem[9][5] ), .B(n6912), .Y(n123) );
  OAI21X1 U170 ( .A(n6465), .B(n6909), .C(n124), .Y(n2580) );
  NAND2X1 U171 ( .A(\Mem[9][6] ), .B(n6912), .Y(n124) );
  OAI21X1 U172 ( .A(n6460), .B(n6909), .C(n125), .Y(n2581) );
  NAND2X1 U173 ( .A(\Mem[9][7] ), .B(n6912), .Y(n125) );
  OAI21X1 U174 ( .A(n6455), .B(n6909), .C(n126), .Y(n2582) );
  NAND2X1 U175 ( .A(\Mem[9][8] ), .B(n6912), .Y(n126) );
  OAI21X1 U176 ( .A(n6450), .B(n6909), .C(n127), .Y(n2583) );
  NAND2X1 U177 ( .A(\Mem[9][9] ), .B(n6912), .Y(n127) );
  OAI21X1 U178 ( .A(n6600), .B(n6909), .C(n128), .Y(n2584) );
  NAND2X1 U179 ( .A(\Mem[9][10] ), .B(n6912), .Y(n128) );
  OAI21X1 U180 ( .A(n6595), .B(n6909), .C(n129), .Y(n2585) );
  NAND2X1 U181 ( .A(\Mem[9][11] ), .B(n6912), .Y(n129) );
  OAI21X1 U182 ( .A(n6590), .B(n6909), .C(n130), .Y(n2586) );
  NAND2X1 U183 ( .A(\Mem[9][12] ), .B(n6912), .Y(n130) );
  OAI21X1 U184 ( .A(n6585), .B(n6910), .C(n131), .Y(n2587) );
  NAND2X1 U185 ( .A(\Mem[9][13] ), .B(n6912), .Y(n131) );
  OAI21X1 U186 ( .A(n6580), .B(n6910), .C(n132), .Y(n2588) );
  NAND2X1 U187 ( .A(\Mem[9][14] ), .B(n6912), .Y(n132) );
  OAI21X1 U188 ( .A(n6575), .B(n6910), .C(n133), .Y(n2589) );
  NAND2X1 U189 ( .A(\Mem[9][15] ), .B(n6911), .Y(n133) );
  OAI21X1 U190 ( .A(n6570), .B(n6910), .C(n134), .Y(n2590) );
  NAND2X1 U191 ( .A(\Mem[9][16] ), .B(n6912), .Y(n134) );
  OAI21X1 U192 ( .A(n6565), .B(n6910), .C(n135), .Y(n2591) );
  NAND2X1 U193 ( .A(\Mem[9][17] ), .B(n6911), .Y(n135) );
  OAI21X1 U194 ( .A(n6560), .B(n6910), .C(n136), .Y(n2592) );
  NAND2X1 U195 ( .A(\Mem[9][18] ), .B(n6911), .Y(n136) );
  OAI21X1 U196 ( .A(n6554), .B(n6910), .C(n137), .Y(n2593) );
  NAND2X1 U197 ( .A(\Mem[9][19] ), .B(n6911), .Y(n137) );
  OAI21X1 U198 ( .A(n6544), .B(n6910), .C(n138), .Y(n2594) );
  NAND2X1 U199 ( .A(\Mem[9][20] ), .B(n6911), .Y(n138) );
  OAI21X1 U200 ( .A(n6539), .B(n6910), .C(n139), .Y(n2595) );
  NAND2X1 U201 ( .A(\Mem[9][21] ), .B(n6911), .Y(n139) );
  OAI21X1 U202 ( .A(n6534), .B(n6910), .C(n140), .Y(n2596) );
  NAND2X1 U203 ( .A(\Mem[9][22] ), .B(n6912), .Y(n140) );
  OAI21X1 U204 ( .A(n6529), .B(n6911), .C(n141), .Y(n2597) );
  NAND2X1 U205 ( .A(\Mem[9][23] ), .B(n6911), .Y(n141) );
  OAI21X1 U206 ( .A(n6524), .B(n6910), .C(n142), .Y(n2598) );
  NAND2X1 U207 ( .A(\Mem[9][24] ), .B(n6912), .Y(n142) );
  OAI21X1 U208 ( .A(n6519), .B(n6911), .C(n143), .Y(n2599) );
  NAND2X1 U209 ( .A(\Mem[9][25] ), .B(n6912), .Y(n143) );
  OAI21X1 U210 ( .A(n6514), .B(n6911), .C(n144), .Y(n2600) );
  NAND2X1 U211 ( .A(\Mem[9][26] ), .B(n6912), .Y(n144) );
  OAI21X1 U212 ( .A(n6509), .B(n6911), .C(n145), .Y(n2601) );
  NAND2X1 U213 ( .A(\Mem[9][27] ), .B(n6912), .Y(n145) );
  OAI21X1 U214 ( .A(n6504), .B(n6911), .C(n146), .Y(n2602) );
  NAND2X1 U215 ( .A(\Mem[9][28] ), .B(n6912), .Y(n146) );
  OAI21X1 U216 ( .A(n6499), .B(n6911), .C(n147), .Y(n2603) );
  NAND2X1 U217 ( .A(\Mem[9][29] ), .B(n6912), .Y(n147) );
  OAI21X1 U218 ( .A(n6489), .B(n6911), .C(n148), .Y(n2604) );
  NAND2X1 U219 ( .A(\Mem[9][30] ), .B(n6913), .Y(n148) );
  OAI21X1 U220 ( .A(n6484), .B(n6911), .C(n149), .Y(n2605) );
  NAND2X1 U221 ( .A(\Mem[9][31] ), .B(n6913), .Y(n149) );
  NAND2X1 U222 ( .A(n7017), .B(n7007), .Y(n117) );
  OAI21X1 U223 ( .A(n6604), .B(n6905), .C(n152), .Y(n2606) );
  NAND2X1 U224 ( .A(\Mem[10][0] ), .B(n6908), .Y(n152) );
  OAI21X1 U225 ( .A(n6549), .B(n6904), .C(n153), .Y(n2607) );
  NAND2X1 U226 ( .A(\Mem[10][1] ), .B(n6908), .Y(n153) );
  OAI21X1 U227 ( .A(n6494), .B(n6904), .C(n154), .Y(n2608) );
  NAND2X1 U228 ( .A(\Mem[10][2] ), .B(n6908), .Y(n154) );
  OAI21X1 U229 ( .A(n6479), .B(n6904), .C(n155), .Y(n2609) );
  NAND2X1 U230 ( .A(\Mem[10][3] ), .B(n6907), .Y(n155) );
  OAI21X1 U231 ( .A(n6474), .B(n6904), .C(n156), .Y(n2610) );
  NAND2X1 U232 ( .A(\Mem[10][4] ), .B(n6908), .Y(n156) );
  OAI21X1 U233 ( .A(n6469), .B(n6904), .C(n157), .Y(n2611) );
  NAND2X1 U234 ( .A(\Mem[10][5] ), .B(n6907), .Y(n157) );
  OAI21X1 U235 ( .A(n6464), .B(n6904), .C(n158), .Y(n2612) );
  NAND2X1 U236 ( .A(\Mem[10][6] ), .B(n6907), .Y(n158) );
  OAI21X1 U237 ( .A(n6459), .B(n6904), .C(n159), .Y(n2613) );
  NAND2X1 U238 ( .A(\Mem[10][7] ), .B(n6907), .Y(n159) );
  OAI21X1 U239 ( .A(n6454), .B(n6904), .C(n160), .Y(n2614) );
  NAND2X1 U240 ( .A(\Mem[10][8] ), .B(n6907), .Y(n160) );
  OAI21X1 U241 ( .A(n6449), .B(n6904), .C(n161), .Y(n2615) );
  NAND2X1 U242 ( .A(\Mem[10][9] ), .B(n6907), .Y(n161) );
  OAI21X1 U243 ( .A(n6599), .B(n6904), .C(n162), .Y(n2616) );
  NAND2X1 U244 ( .A(\Mem[10][10] ), .B(n6907), .Y(n162) );
  OAI21X1 U245 ( .A(n6594), .B(n6904), .C(n163), .Y(n2617) );
  NAND2X1 U246 ( .A(\Mem[10][11] ), .B(n6907), .Y(n163) );
  OAI21X1 U247 ( .A(n6589), .B(n6904), .C(n164), .Y(n2618) );
  NAND2X1 U248 ( .A(\Mem[10][12] ), .B(n6907), .Y(n164) );
  OAI21X1 U249 ( .A(n6584), .B(n6905), .C(n165), .Y(n2619) );
  NAND2X1 U250 ( .A(\Mem[10][13] ), .B(n6907), .Y(n165) );
  OAI21X1 U251 ( .A(n6579), .B(n6905), .C(n166), .Y(n2620) );
  NAND2X1 U252 ( .A(\Mem[10][14] ), .B(n6907), .Y(n166) );
  OAI21X1 U253 ( .A(n6574), .B(n6905), .C(n167), .Y(n2621) );
  NAND2X1 U254 ( .A(\Mem[10][15] ), .B(n6906), .Y(n167) );
  OAI21X1 U255 ( .A(n6569), .B(n6905), .C(n168), .Y(n2622) );
  NAND2X1 U256 ( .A(\Mem[10][16] ), .B(n6907), .Y(n168) );
  OAI21X1 U257 ( .A(n6564), .B(n6905), .C(n169), .Y(n2623) );
  NAND2X1 U258 ( .A(\Mem[10][17] ), .B(n6906), .Y(n169) );
  OAI21X1 U259 ( .A(n6559), .B(n6905), .C(n170), .Y(n2624) );
  NAND2X1 U260 ( .A(\Mem[10][18] ), .B(n6906), .Y(n170) );
  OAI21X1 U261 ( .A(n6554), .B(n6905), .C(n171), .Y(n2625) );
  NAND2X1 U262 ( .A(\Mem[10][19] ), .B(n6906), .Y(n171) );
  OAI21X1 U263 ( .A(n6544), .B(n6905), .C(n172), .Y(n2626) );
  NAND2X1 U264 ( .A(\Mem[10][20] ), .B(n6906), .Y(n172) );
  OAI21X1 U265 ( .A(n6539), .B(n6905), .C(n173), .Y(n2627) );
  NAND2X1 U266 ( .A(\Mem[10][21] ), .B(n6906), .Y(n173) );
  OAI21X1 U267 ( .A(n6534), .B(n6905), .C(n174), .Y(n2628) );
  NAND2X1 U268 ( .A(\Mem[10][22] ), .B(n6907), .Y(n174) );
  OAI21X1 U269 ( .A(n6529), .B(n6906), .C(n175), .Y(n2629) );
  NAND2X1 U270 ( .A(\Mem[10][23] ), .B(n6906), .Y(n175) );
  OAI21X1 U271 ( .A(n6524), .B(n6905), .C(n176), .Y(n2630) );
  NAND2X1 U272 ( .A(\Mem[10][24] ), .B(n6907), .Y(n176) );
  OAI21X1 U273 ( .A(n6519), .B(n6906), .C(n177), .Y(n2631) );
  NAND2X1 U274 ( .A(\Mem[10][25] ), .B(n6907), .Y(n177) );
  OAI21X1 U275 ( .A(n6514), .B(n6906), .C(n178), .Y(n2632) );
  NAND2X1 U276 ( .A(\Mem[10][26] ), .B(n6907), .Y(n178) );
  OAI21X1 U277 ( .A(n6509), .B(n6906), .C(n179), .Y(n2633) );
  NAND2X1 U278 ( .A(\Mem[10][27] ), .B(n6907), .Y(n179) );
  OAI21X1 U279 ( .A(n6504), .B(n6906), .C(n180), .Y(n2634) );
  NAND2X1 U280 ( .A(\Mem[10][28] ), .B(n6907), .Y(n180) );
  OAI21X1 U281 ( .A(n6499), .B(n6906), .C(n181), .Y(n2635) );
  NAND2X1 U282 ( .A(\Mem[10][29] ), .B(n6907), .Y(n181) );
  OAI21X1 U283 ( .A(n6489), .B(n6906), .C(n182), .Y(n2636) );
  NAND2X1 U284 ( .A(\Mem[10][30] ), .B(n6908), .Y(n182) );
  OAI21X1 U285 ( .A(n6484), .B(n6906), .C(n183), .Y(n2637) );
  NAND2X1 U286 ( .A(\Mem[10][31] ), .B(n6908), .Y(n183) );
  NAND2X1 U287 ( .A(n7018), .B(n7007), .Y(n151) );
  OAI21X1 U288 ( .A(n6604), .B(n6900), .C(n186), .Y(n2638) );
  NAND2X1 U289 ( .A(\Mem[11][0] ), .B(n6903), .Y(n186) );
  OAI21X1 U290 ( .A(n6549), .B(n6899), .C(n187), .Y(n2639) );
  NAND2X1 U291 ( .A(\Mem[11][1] ), .B(n6903), .Y(n187) );
  OAI21X1 U292 ( .A(n6494), .B(n6899), .C(n188), .Y(n2640) );
  NAND2X1 U293 ( .A(\Mem[11][2] ), .B(n6903), .Y(n188) );
  OAI21X1 U294 ( .A(n6479), .B(n6899), .C(n189), .Y(n2641) );
  NAND2X1 U295 ( .A(\Mem[11][3] ), .B(n6902), .Y(n189) );
  OAI21X1 U296 ( .A(n6474), .B(n6899), .C(n190), .Y(n2642) );
  NAND2X1 U297 ( .A(\Mem[11][4] ), .B(n6903), .Y(n190) );
  OAI21X1 U298 ( .A(n6469), .B(n6899), .C(n191), .Y(n2643) );
  NAND2X1 U299 ( .A(\Mem[11][5] ), .B(n6902), .Y(n191) );
  OAI21X1 U300 ( .A(n6464), .B(n6899), .C(n192), .Y(n2644) );
  NAND2X1 U301 ( .A(\Mem[11][6] ), .B(n6902), .Y(n192) );
  OAI21X1 U302 ( .A(n6459), .B(n6899), .C(n193), .Y(n2645) );
  NAND2X1 U303 ( .A(\Mem[11][7] ), .B(n6902), .Y(n193) );
  OAI21X1 U304 ( .A(n6454), .B(n6899), .C(n194), .Y(n2646) );
  NAND2X1 U305 ( .A(\Mem[11][8] ), .B(n6902), .Y(n194) );
  OAI21X1 U306 ( .A(n6449), .B(n6899), .C(n195), .Y(n2647) );
  NAND2X1 U307 ( .A(\Mem[11][9] ), .B(n6902), .Y(n195) );
  OAI21X1 U308 ( .A(n6599), .B(n6899), .C(n196), .Y(n2648) );
  NAND2X1 U309 ( .A(\Mem[11][10] ), .B(n6902), .Y(n196) );
  OAI21X1 U310 ( .A(n6594), .B(n6899), .C(n197), .Y(n2649) );
  NAND2X1 U311 ( .A(\Mem[11][11] ), .B(n6902), .Y(n197) );
  OAI21X1 U312 ( .A(n6589), .B(n6899), .C(n198), .Y(n2650) );
  NAND2X1 U313 ( .A(\Mem[11][12] ), .B(n6902), .Y(n198) );
  OAI21X1 U314 ( .A(n6584), .B(n6900), .C(n199), .Y(n2651) );
  NAND2X1 U315 ( .A(\Mem[11][13] ), .B(n6902), .Y(n199) );
  OAI21X1 U316 ( .A(n6579), .B(n6900), .C(n200), .Y(n2652) );
  NAND2X1 U317 ( .A(\Mem[11][14] ), .B(n6902), .Y(n200) );
  OAI21X1 U318 ( .A(n6574), .B(n6900), .C(n201), .Y(n2653) );
  NAND2X1 U319 ( .A(\Mem[11][15] ), .B(n6901), .Y(n201) );
  OAI21X1 U320 ( .A(n6569), .B(n6900), .C(n202), .Y(n2654) );
  NAND2X1 U321 ( .A(\Mem[11][16] ), .B(n6902), .Y(n202) );
  OAI21X1 U322 ( .A(n6564), .B(n6900), .C(n203), .Y(n2655) );
  NAND2X1 U323 ( .A(\Mem[11][17] ), .B(n6901), .Y(n203) );
  OAI21X1 U324 ( .A(n6559), .B(n6900), .C(n204), .Y(n2656) );
  NAND2X1 U325 ( .A(\Mem[11][18] ), .B(n6901), .Y(n204) );
  OAI21X1 U326 ( .A(n6554), .B(n6900), .C(n205), .Y(n2657) );
  NAND2X1 U327 ( .A(\Mem[11][19] ), .B(n6901), .Y(n205) );
  OAI21X1 U328 ( .A(n6544), .B(n6900), .C(n206), .Y(n2658) );
  NAND2X1 U329 ( .A(\Mem[11][20] ), .B(n6901), .Y(n206) );
  OAI21X1 U330 ( .A(n6539), .B(n6900), .C(n207), .Y(n2659) );
  NAND2X1 U331 ( .A(\Mem[11][21] ), .B(n6901), .Y(n207) );
  OAI21X1 U332 ( .A(n6534), .B(n6900), .C(n208), .Y(n2660) );
  NAND2X1 U333 ( .A(\Mem[11][22] ), .B(n6902), .Y(n208) );
  OAI21X1 U334 ( .A(n6529), .B(n6901), .C(n209), .Y(n2661) );
  NAND2X1 U335 ( .A(\Mem[11][23] ), .B(n6901), .Y(n209) );
  OAI21X1 U336 ( .A(n6524), .B(n6900), .C(n210), .Y(n2662) );
  NAND2X1 U337 ( .A(\Mem[11][24] ), .B(n6902), .Y(n210) );
  OAI21X1 U338 ( .A(n6519), .B(n6901), .C(n211), .Y(n2663) );
  NAND2X1 U339 ( .A(\Mem[11][25] ), .B(n6902), .Y(n211) );
  OAI21X1 U340 ( .A(n6514), .B(n6901), .C(n212), .Y(n2664) );
  NAND2X1 U341 ( .A(\Mem[11][26] ), .B(n6902), .Y(n212) );
  OAI21X1 U342 ( .A(n6509), .B(n6901), .C(n213), .Y(n2665) );
  NAND2X1 U343 ( .A(\Mem[11][27] ), .B(n6902), .Y(n213) );
  OAI21X1 U344 ( .A(n6504), .B(n6901), .C(n214), .Y(n2666) );
  NAND2X1 U345 ( .A(\Mem[11][28] ), .B(n6902), .Y(n214) );
  OAI21X1 U346 ( .A(n6499), .B(n6901), .C(n215), .Y(n2667) );
  NAND2X1 U347 ( .A(\Mem[11][29] ), .B(n6902), .Y(n215) );
  OAI21X1 U348 ( .A(n6489), .B(n6901), .C(n216), .Y(n2668) );
  NAND2X1 U349 ( .A(\Mem[11][30] ), .B(n6903), .Y(n216) );
  OAI21X1 U350 ( .A(n6484), .B(n6901), .C(n217), .Y(n2669) );
  NAND2X1 U351 ( .A(\Mem[11][31] ), .B(n6903), .Y(n217) );
  NAND2X1 U352 ( .A(n7019), .B(n7007), .Y(n185) );
  OAI21X1 U353 ( .A(n6604), .B(n6895), .C(n220), .Y(n2670) );
  NAND2X1 U354 ( .A(\Mem[12][0] ), .B(n6898), .Y(n220) );
  OAI21X1 U355 ( .A(n6549), .B(n6894), .C(n221), .Y(n2671) );
  NAND2X1 U356 ( .A(\Mem[12][1] ), .B(n6898), .Y(n221) );
  OAI21X1 U357 ( .A(n6494), .B(n6894), .C(n222), .Y(n2672) );
  NAND2X1 U358 ( .A(\Mem[12][2] ), .B(n6898), .Y(n222) );
  OAI21X1 U359 ( .A(n6479), .B(n6894), .C(n223), .Y(n2673) );
  NAND2X1 U360 ( .A(\Mem[12][3] ), .B(n6897), .Y(n223) );
  OAI21X1 U361 ( .A(n6474), .B(n6894), .C(n224), .Y(n2674) );
  NAND2X1 U362 ( .A(\Mem[12][4] ), .B(n6898), .Y(n224) );
  OAI21X1 U363 ( .A(n6469), .B(n6894), .C(n225), .Y(n2675) );
  NAND2X1 U364 ( .A(\Mem[12][5] ), .B(n6897), .Y(n225) );
  OAI21X1 U365 ( .A(n6464), .B(n6894), .C(n226), .Y(n2676) );
  NAND2X1 U366 ( .A(\Mem[12][6] ), .B(n6897), .Y(n226) );
  OAI21X1 U367 ( .A(n6459), .B(n6894), .C(n227), .Y(n2677) );
  NAND2X1 U368 ( .A(\Mem[12][7] ), .B(n6897), .Y(n227) );
  OAI21X1 U369 ( .A(n6454), .B(n6894), .C(n228), .Y(n2678) );
  NAND2X1 U370 ( .A(\Mem[12][8] ), .B(n6897), .Y(n228) );
  OAI21X1 U371 ( .A(n6449), .B(n6894), .C(n229), .Y(n2679) );
  NAND2X1 U372 ( .A(\Mem[12][9] ), .B(n6897), .Y(n229) );
  OAI21X1 U373 ( .A(n6599), .B(n6894), .C(n230), .Y(n2680) );
  NAND2X1 U374 ( .A(\Mem[12][10] ), .B(n6897), .Y(n230) );
  OAI21X1 U375 ( .A(n6594), .B(n6894), .C(n231), .Y(n2681) );
  NAND2X1 U376 ( .A(\Mem[12][11] ), .B(n6897), .Y(n231) );
  OAI21X1 U377 ( .A(n6589), .B(n6894), .C(n232), .Y(n2682) );
  NAND2X1 U378 ( .A(\Mem[12][12] ), .B(n6897), .Y(n232) );
  OAI21X1 U379 ( .A(n6584), .B(n6895), .C(n233), .Y(n2683) );
  NAND2X1 U380 ( .A(\Mem[12][13] ), .B(n6897), .Y(n233) );
  OAI21X1 U381 ( .A(n6579), .B(n6895), .C(n234), .Y(n2684) );
  NAND2X1 U382 ( .A(\Mem[12][14] ), .B(n6897), .Y(n234) );
  OAI21X1 U383 ( .A(n6574), .B(n6895), .C(n235), .Y(n2685) );
  NAND2X1 U384 ( .A(\Mem[12][15] ), .B(n6896), .Y(n235) );
  OAI21X1 U385 ( .A(n6569), .B(n6895), .C(n236), .Y(n2686) );
  NAND2X1 U386 ( .A(\Mem[12][16] ), .B(n6897), .Y(n236) );
  OAI21X1 U387 ( .A(n6564), .B(n6895), .C(n237), .Y(n2687) );
  NAND2X1 U388 ( .A(\Mem[12][17] ), .B(n6896), .Y(n237) );
  OAI21X1 U389 ( .A(n6559), .B(n6895), .C(n238), .Y(n2688) );
  NAND2X1 U390 ( .A(\Mem[12][18] ), .B(n6896), .Y(n238) );
  OAI21X1 U391 ( .A(n6554), .B(n6895), .C(n239), .Y(n2689) );
  NAND2X1 U392 ( .A(\Mem[12][19] ), .B(n6896), .Y(n239) );
  OAI21X1 U393 ( .A(n6544), .B(n6895), .C(n240), .Y(n2690) );
  NAND2X1 U394 ( .A(\Mem[12][20] ), .B(n6896), .Y(n240) );
  OAI21X1 U395 ( .A(n6539), .B(n6895), .C(n241), .Y(n2691) );
  NAND2X1 U396 ( .A(\Mem[12][21] ), .B(n6896), .Y(n241) );
  OAI21X1 U397 ( .A(n6534), .B(n6895), .C(n242), .Y(n2692) );
  NAND2X1 U398 ( .A(\Mem[12][22] ), .B(n6897), .Y(n242) );
  OAI21X1 U399 ( .A(n6529), .B(n6896), .C(n243), .Y(n2693) );
  NAND2X1 U400 ( .A(\Mem[12][23] ), .B(n6896), .Y(n243) );
  OAI21X1 U401 ( .A(n6524), .B(n6895), .C(n244), .Y(n2694) );
  NAND2X1 U402 ( .A(\Mem[12][24] ), .B(n6897), .Y(n244) );
  OAI21X1 U403 ( .A(n6519), .B(n6896), .C(n245), .Y(n2695) );
  NAND2X1 U404 ( .A(\Mem[12][25] ), .B(n6897), .Y(n245) );
  OAI21X1 U405 ( .A(n6514), .B(n6896), .C(n246), .Y(n2696) );
  NAND2X1 U406 ( .A(\Mem[12][26] ), .B(n6897), .Y(n246) );
  OAI21X1 U407 ( .A(n6509), .B(n6896), .C(n247), .Y(n2697) );
  NAND2X1 U408 ( .A(\Mem[12][27] ), .B(n6897), .Y(n247) );
  OAI21X1 U409 ( .A(n6504), .B(n6896), .C(n248), .Y(n2698) );
  NAND2X1 U410 ( .A(\Mem[12][28] ), .B(n6897), .Y(n248) );
  OAI21X1 U411 ( .A(n6499), .B(n6896), .C(n249), .Y(n2699) );
  NAND2X1 U412 ( .A(\Mem[12][29] ), .B(n6897), .Y(n249) );
  OAI21X1 U413 ( .A(n6489), .B(n6896), .C(n250), .Y(n2700) );
  NAND2X1 U414 ( .A(\Mem[12][30] ), .B(n6898), .Y(n250) );
  OAI21X1 U415 ( .A(n6484), .B(n6896), .C(n251), .Y(n2701) );
  NAND2X1 U416 ( .A(\Mem[12][31] ), .B(n6898), .Y(n251) );
  NAND2X1 U417 ( .A(n7022), .B(n7007), .Y(n219) );
  OAI21X1 U418 ( .A(n6604), .B(n6890), .C(n254), .Y(n2702) );
  NAND2X1 U419 ( .A(\Mem[13][0] ), .B(n6893), .Y(n254) );
  OAI21X1 U420 ( .A(n6549), .B(n6889), .C(n255), .Y(n2703) );
  NAND2X1 U421 ( .A(\Mem[13][1] ), .B(n6893), .Y(n255) );
  OAI21X1 U422 ( .A(n6494), .B(n6889), .C(n256), .Y(n2704) );
  NAND2X1 U423 ( .A(\Mem[13][2] ), .B(n6893), .Y(n256) );
  OAI21X1 U424 ( .A(n6479), .B(n6889), .C(n257), .Y(n2705) );
  NAND2X1 U425 ( .A(\Mem[13][3] ), .B(n6892), .Y(n257) );
  OAI21X1 U426 ( .A(n6474), .B(n6889), .C(n258), .Y(n2706) );
  NAND2X1 U427 ( .A(\Mem[13][4] ), .B(n6893), .Y(n258) );
  OAI21X1 U428 ( .A(n6469), .B(n6889), .C(n259), .Y(n2707) );
  NAND2X1 U429 ( .A(\Mem[13][5] ), .B(n6892), .Y(n259) );
  OAI21X1 U430 ( .A(n6464), .B(n6889), .C(n260), .Y(n2708) );
  NAND2X1 U431 ( .A(\Mem[13][6] ), .B(n6892), .Y(n260) );
  OAI21X1 U432 ( .A(n6459), .B(n6889), .C(n261), .Y(n2709) );
  NAND2X1 U433 ( .A(\Mem[13][7] ), .B(n6892), .Y(n261) );
  OAI21X1 U434 ( .A(n6454), .B(n6889), .C(n262), .Y(n2710) );
  NAND2X1 U435 ( .A(\Mem[13][8] ), .B(n6892), .Y(n262) );
  OAI21X1 U436 ( .A(n6449), .B(n6889), .C(n263), .Y(n2711) );
  NAND2X1 U437 ( .A(\Mem[13][9] ), .B(n6892), .Y(n263) );
  OAI21X1 U438 ( .A(n6599), .B(n6889), .C(n264), .Y(n2712) );
  NAND2X1 U439 ( .A(\Mem[13][10] ), .B(n6892), .Y(n264) );
  OAI21X1 U440 ( .A(n6594), .B(n6889), .C(n265), .Y(n2713) );
  NAND2X1 U441 ( .A(\Mem[13][11] ), .B(n6892), .Y(n265) );
  OAI21X1 U442 ( .A(n6589), .B(n6889), .C(n266), .Y(n2714) );
  NAND2X1 U443 ( .A(\Mem[13][12] ), .B(n6892), .Y(n266) );
  OAI21X1 U444 ( .A(n6584), .B(n6890), .C(n267), .Y(n2715) );
  NAND2X1 U445 ( .A(\Mem[13][13] ), .B(n6892), .Y(n267) );
  OAI21X1 U446 ( .A(n6579), .B(n6890), .C(n268), .Y(n2716) );
  NAND2X1 U447 ( .A(\Mem[13][14] ), .B(n6892), .Y(n268) );
  OAI21X1 U448 ( .A(n6574), .B(n6890), .C(n269), .Y(n2717) );
  NAND2X1 U449 ( .A(\Mem[13][15] ), .B(n6891), .Y(n269) );
  OAI21X1 U450 ( .A(n6569), .B(n6890), .C(n270), .Y(n2718) );
  NAND2X1 U451 ( .A(\Mem[13][16] ), .B(n6892), .Y(n270) );
  OAI21X1 U452 ( .A(n6564), .B(n6890), .C(n271), .Y(n2719) );
  NAND2X1 U453 ( .A(\Mem[13][17] ), .B(n6891), .Y(n271) );
  OAI21X1 U454 ( .A(n6559), .B(n6890), .C(n272), .Y(n2720) );
  NAND2X1 U455 ( .A(\Mem[13][18] ), .B(n6891), .Y(n272) );
  OAI21X1 U456 ( .A(n6554), .B(n6890), .C(n273), .Y(n2721) );
  NAND2X1 U457 ( .A(\Mem[13][19] ), .B(n6891), .Y(n273) );
  OAI21X1 U458 ( .A(n6544), .B(n6890), .C(n274), .Y(n2722) );
  NAND2X1 U459 ( .A(\Mem[13][20] ), .B(n6891), .Y(n274) );
  OAI21X1 U460 ( .A(n6539), .B(n6890), .C(n275), .Y(n2723) );
  NAND2X1 U461 ( .A(\Mem[13][21] ), .B(n6891), .Y(n275) );
  OAI21X1 U462 ( .A(n6534), .B(n6890), .C(n276), .Y(n2724) );
  NAND2X1 U463 ( .A(\Mem[13][22] ), .B(n6892), .Y(n276) );
  OAI21X1 U464 ( .A(n6529), .B(n6891), .C(n277), .Y(n2725) );
  NAND2X1 U465 ( .A(\Mem[13][23] ), .B(n6891), .Y(n277) );
  OAI21X1 U466 ( .A(n6524), .B(n6890), .C(n278), .Y(n2726) );
  NAND2X1 U467 ( .A(\Mem[13][24] ), .B(n6892), .Y(n278) );
  OAI21X1 U468 ( .A(n6519), .B(n6891), .C(n279), .Y(n2727) );
  NAND2X1 U469 ( .A(\Mem[13][25] ), .B(n6892), .Y(n279) );
  OAI21X1 U470 ( .A(n6514), .B(n6891), .C(n280), .Y(n2728) );
  NAND2X1 U471 ( .A(\Mem[13][26] ), .B(n6892), .Y(n280) );
  OAI21X1 U472 ( .A(n6509), .B(n6891), .C(n281), .Y(n2729) );
  NAND2X1 U473 ( .A(\Mem[13][27] ), .B(n6892), .Y(n281) );
  OAI21X1 U474 ( .A(n6504), .B(n6891), .C(n282), .Y(n2730) );
  NAND2X1 U475 ( .A(\Mem[13][28] ), .B(n6892), .Y(n282) );
  OAI21X1 U476 ( .A(n6499), .B(n6891), .C(n283), .Y(n2731) );
  NAND2X1 U477 ( .A(\Mem[13][29] ), .B(n6892), .Y(n283) );
  OAI21X1 U478 ( .A(n6489), .B(n6891), .C(n284), .Y(n2732) );
  NAND2X1 U479 ( .A(\Mem[13][30] ), .B(n6893), .Y(n284) );
  OAI21X1 U480 ( .A(n6484), .B(n6891), .C(n285), .Y(n2733) );
  NAND2X1 U481 ( .A(\Mem[13][31] ), .B(n6893), .Y(n285) );
  NAND2X1 U482 ( .A(n7023), .B(n7007), .Y(n253) );
  OAI21X1 U483 ( .A(n6604), .B(n6885), .C(n288), .Y(n2734) );
  NAND2X1 U484 ( .A(\Mem[14][0] ), .B(n6888), .Y(n288) );
  OAI21X1 U485 ( .A(n6549), .B(n6884), .C(n289), .Y(n2735) );
  NAND2X1 U486 ( .A(\Mem[14][1] ), .B(n6888), .Y(n289) );
  OAI21X1 U487 ( .A(n6494), .B(n6884), .C(n290), .Y(n2736) );
  NAND2X1 U488 ( .A(\Mem[14][2] ), .B(n6888), .Y(n290) );
  OAI21X1 U489 ( .A(n6479), .B(n6884), .C(n291), .Y(n2737) );
  NAND2X1 U490 ( .A(\Mem[14][3] ), .B(n6887), .Y(n291) );
  OAI21X1 U491 ( .A(n6474), .B(n6884), .C(n292), .Y(n2738) );
  NAND2X1 U492 ( .A(\Mem[14][4] ), .B(n6888), .Y(n292) );
  OAI21X1 U493 ( .A(n6469), .B(n6884), .C(n293), .Y(n2739) );
  NAND2X1 U494 ( .A(\Mem[14][5] ), .B(n6887), .Y(n293) );
  OAI21X1 U495 ( .A(n6464), .B(n6884), .C(n294), .Y(n2740) );
  NAND2X1 U496 ( .A(\Mem[14][6] ), .B(n6887), .Y(n294) );
  OAI21X1 U497 ( .A(n6459), .B(n6884), .C(n295), .Y(n2741) );
  NAND2X1 U498 ( .A(\Mem[14][7] ), .B(n6887), .Y(n295) );
  OAI21X1 U499 ( .A(n6454), .B(n6884), .C(n296), .Y(n2742) );
  NAND2X1 U500 ( .A(\Mem[14][8] ), .B(n6887), .Y(n296) );
  OAI21X1 U501 ( .A(n6449), .B(n6884), .C(n297), .Y(n2743) );
  NAND2X1 U502 ( .A(\Mem[14][9] ), .B(n6887), .Y(n297) );
  OAI21X1 U503 ( .A(n6599), .B(n6884), .C(n298), .Y(n2744) );
  NAND2X1 U504 ( .A(\Mem[14][10] ), .B(n6887), .Y(n298) );
  OAI21X1 U505 ( .A(n6594), .B(n6884), .C(n299), .Y(n2745) );
  NAND2X1 U506 ( .A(\Mem[14][11] ), .B(n6887), .Y(n299) );
  OAI21X1 U507 ( .A(n6589), .B(n6884), .C(n300), .Y(n2746) );
  NAND2X1 U508 ( .A(\Mem[14][12] ), .B(n6887), .Y(n300) );
  OAI21X1 U509 ( .A(n6584), .B(n6885), .C(n301), .Y(n2747) );
  NAND2X1 U510 ( .A(\Mem[14][13] ), .B(n6887), .Y(n301) );
  OAI21X1 U511 ( .A(n6579), .B(n6885), .C(n302), .Y(n2748) );
  NAND2X1 U512 ( .A(\Mem[14][14] ), .B(n6887), .Y(n302) );
  OAI21X1 U513 ( .A(n6574), .B(n6885), .C(n303), .Y(n2749) );
  NAND2X1 U514 ( .A(\Mem[14][15] ), .B(n6886), .Y(n303) );
  OAI21X1 U515 ( .A(n6569), .B(n6885), .C(n304), .Y(n2750) );
  NAND2X1 U516 ( .A(\Mem[14][16] ), .B(n6887), .Y(n304) );
  OAI21X1 U517 ( .A(n6564), .B(n6885), .C(n305), .Y(n2751) );
  NAND2X1 U518 ( .A(\Mem[14][17] ), .B(n6886), .Y(n305) );
  OAI21X1 U519 ( .A(n6559), .B(n6885), .C(n306), .Y(n2752) );
  NAND2X1 U520 ( .A(\Mem[14][18] ), .B(n6886), .Y(n306) );
  OAI21X1 U521 ( .A(n6554), .B(n6885), .C(n307), .Y(n2753) );
  NAND2X1 U522 ( .A(\Mem[14][19] ), .B(n6886), .Y(n307) );
  OAI21X1 U523 ( .A(n6544), .B(n6885), .C(n308), .Y(n2754) );
  NAND2X1 U524 ( .A(\Mem[14][20] ), .B(n6886), .Y(n308) );
  OAI21X1 U525 ( .A(n6539), .B(n6885), .C(n309), .Y(n2755) );
  NAND2X1 U526 ( .A(\Mem[14][21] ), .B(n6886), .Y(n309) );
  OAI21X1 U527 ( .A(n6534), .B(n6885), .C(n310), .Y(n2756) );
  NAND2X1 U528 ( .A(\Mem[14][22] ), .B(n6887), .Y(n310) );
  OAI21X1 U529 ( .A(n6529), .B(n6886), .C(n311), .Y(n2757) );
  NAND2X1 U530 ( .A(\Mem[14][23] ), .B(n6886), .Y(n311) );
  OAI21X1 U531 ( .A(n6524), .B(n6885), .C(n312), .Y(n2758) );
  NAND2X1 U532 ( .A(\Mem[14][24] ), .B(n6887), .Y(n312) );
  OAI21X1 U533 ( .A(n6519), .B(n6886), .C(n313), .Y(n2759) );
  NAND2X1 U534 ( .A(\Mem[14][25] ), .B(n6887), .Y(n313) );
  OAI21X1 U535 ( .A(n6514), .B(n6886), .C(n314), .Y(n2760) );
  NAND2X1 U536 ( .A(\Mem[14][26] ), .B(n6887), .Y(n314) );
  OAI21X1 U537 ( .A(n6509), .B(n6886), .C(n315), .Y(n2761) );
  NAND2X1 U538 ( .A(\Mem[14][27] ), .B(n6887), .Y(n315) );
  OAI21X1 U539 ( .A(n6504), .B(n6886), .C(n316), .Y(n2762) );
  NAND2X1 U540 ( .A(\Mem[14][28] ), .B(n6887), .Y(n316) );
  OAI21X1 U541 ( .A(n6499), .B(n6886), .C(n317), .Y(n2763) );
  NAND2X1 U542 ( .A(\Mem[14][29] ), .B(n6887), .Y(n317) );
  OAI21X1 U543 ( .A(n6489), .B(n6886), .C(n318), .Y(n2764) );
  NAND2X1 U544 ( .A(\Mem[14][30] ), .B(n6888), .Y(n318) );
  OAI21X1 U545 ( .A(n6484), .B(n6886), .C(n319), .Y(n2765) );
  NAND2X1 U546 ( .A(\Mem[14][31] ), .B(n6888), .Y(n319) );
  NAND2X1 U547 ( .A(n7007), .B(n7024), .Y(n287) );
  OAI21X1 U548 ( .A(n6604), .B(n6880), .C(n322), .Y(n2766) );
  NAND2X1 U549 ( .A(\Mem[15][0] ), .B(n6883), .Y(n322) );
  OAI21X1 U550 ( .A(n6549), .B(n6879), .C(n323), .Y(n2767) );
  NAND2X1 U551 ( .A(\Mem[15][1] ), .B(n6883), .Y(n323) );
  OAI21X1 U552 ( .A(n6494), .B(n6879), .C(n324), .Y(n2768) );
  NAND2X1 U553 ( .A(\Mem[15][2] ), .B(n6883), .Y(n324) );
  OAI21X1 U554 ( .A(n6479), .B(n6879), .C(n325), .Y(n2769) );
  NAND2X1 U555 ( .A(\Mem[15][3] ), .B(n6882), .Y(n325) );
  OAI21X1 U556 ( .A(n6474), .B(n6879), .C(n326), .Y(n2770) );
  NAND2X1 U557 ( .A(\Mem[15][4] ), .B(n6883), .Y(n326) );
  OAI21X1 U558 ( .A(n6469), .B(n6879), .C(n327), .Y(n2771) );
  NAND2X1 U559 ( .A(\Mem[15][5] ), .B(n6882), .Y(n327) );
  OAI21X1 U560 ( .A(n6464), .B(n6879), .C(n328), .Y(n2772) );
  NAND2X1 U561 ( .A(\Mem[15][6] ), .B(n6882), .Y(n328) );
  OAI21X1 U562 ( .A(n6459), .B(n6879), .C(n329), .Y(n2773) );
  NAND2X1 U563 ( .A(\Mem[15][7] ), .B(n6882), .Y(n329) );
  OAI21X1 U564 ( .A(n6454), .B(n6879), .C(n330), .Y(n2774) );
  NAND2X1 U565 ( .A(\Mem[15][8] ), .B(n6882), .Y(n330) );
  OAI21X1 U566 ( .A(n6449), .B(n6879), .C(n331), .Y(n2775) );
  NAND2X1 U567 ( .A(\Mem[15][9] ), .B(n6882), .Y(n331) );
  OAI21X1 U568 ( .A(n6599), .B(n6879), .C(n332), .Y(n2776) );
  NAND2X1 U569 ( .A(\Mem[15][10] ), .B(n6882), .Y(n332) );
  OAI21X1 U570 ( .A(n6594), .B(n6879), .C(n333), .Y(n2777) );
  NAND2X1 U571 ( .A(\Mem[15][11] ), .B(n6882), .Y(n333) );
  OAI21X1 U572 ( .A(n6589), .B(n6879), .C(n334), .Y(n2778) );
  NAND2X1 U573 ( .A(\Mem[15][12] ), .B(n6882), .Y(n334) );
  OAI21X1 U574 ( .A(n6584), .B(n6880), .C(n335), .Y(n2779) );
  NAND2X1 U575 ( .A(\Mem[15][13] ), .B(n6882), .Y(n335) );
  OAI21X1 U576 ( .A(n6579), .B(n6880), .C(n336), .Y(n2780) );
  NAND2X1 U577 ( .A(\Mem[15][14] ), .B(n6882), .Y(n336) );
  OAI21X1 U578 ( .A(n6574), .B(n6880), .C(n337), .Y(n2781) );
  NAND2X1 U579 ( .A(\Mem[15][15] ), .B(n6881), .Y(n337) );
  OAI21X1 U580 ( .A(n6569), .B(n6880), .C(n338), .Y(n2782) );
  NAND2X1 U581 ( .A(\Mem[15][16] ), .B(n6882), .Y(n338) );
  OAI21X1 U582 ( .A(n6564), .B(n6880), .C(n339), .Y(n2783) );
  NAND2X1 U583 ( .A(\Mem[15][17] ), .B(n6881), .Y(n339) );
  OAI21X1 U584 ( .A(n6559), .B(n6880), .C(n340), .Y(n2784) );
  NAND2X1 U585 ( .A(\Mem[15][18] ), .B(n6881), .Y(n340) );
  OAI21X1 U586 ( .A(n6554), .B(n6880), .C(n341), .Y(n2785) );
  NAND2X1 U587 ( .A(\Mem[15][19] ), .B(n6881), .Y(n341) );
  OAI21X1 U588 ( .A(n6544), .B(n6880), .C(n342), .Y(n2786) );
  NAND2X1 U589 ( .A(\Mem[15][20] ), .B(n6881), .Y(n342) );
  OAI21X1 U590 ( .A(n6539), .B(n6880), .C(n343), .Y(n2787) );
  NAND2X1 U591 ( .A(\Mem[15][21] ), .B(n6881), .Y(n343) );
  OAI21X1 U592 ( .A(n6534), .B(n6880), .C(n344), .Y(n2788) );
  NAND2X1 U593 ( .A(\Mem[15][22] ), .B(n6882), .Y(n344) );
  OAI21X1 U594 ( .A(n6529), .B(n6881), .C(n345), .Y(n2789) );
  NAND2X1 U595 ( .A(\Mem[15][23] ), .B(n6881), .Y(n345) );
  OAI21X1 U596 ( .A(n6524), .B(n6880), .C(n346), .Y(n2790) );
  NAND2X1 U597 ( .A(\Mem[15][24] ), .B(n6882), .Y(n346) );
  OAI21X1 U598 ( .A(n6519), .B(n6881), .C(n347), .Y(n2791) );
  NAND2X1 U599 ( .A(\Mem[15][25] ), .B(n6882), .Y(n347) );
  OAI21X1 U600 ( .A(n6514), .B(n6881), .C(n348), .Y(n2792) );
  NAND2X1 U601 ( .A(\Mem[15][26] ), .B(n6882), .Y(n348) );
  OAI21X1 U602 ( .A(n6509), .B(n6881), .C(n349), .Y(n2793) );
  NAND2X1 U603 ( .A(\Mem[15][27] ), .B(n6882), .Y(n349) );
  OAI21X1 U604 ( .A(n6504), .B(n6881), .C(n350), .Y(n2794) );
  NAND2X1 U605 ( .A(\Mem[15][28] ), .B(n6882), .Y(n350) );
  OAI21X1 U606 ( .A(n6499), .B(n6881), .C(n351), .Y(n2795) );
  NAND2X1 U607 ( .A(\Mem[15][29] ), .B(n6882), .Y(n351) );
  OAI21X1 U608 ( .A(n6489), .B(n6881), .C(n352), .Y(n2796) );
  NAND2X1 U609 ( .A(\Mem[15][30] ), .B(n6883), .Y(n352) );
  OAI21X1 U610 ( .A(n6484), .B(n6881), .C(n353), .Y(n2797) );
  NAND2X1 U611 ( .A(\Mem[15][31] ), .B(n6883), .Y(n353) );
  NAND2X1 U612 ( .A(n7007), .B(n7021), .Y(n321) );
  NAND3X1 U614 ( .A(n355), .B(n7014), .C(ADDR_WR[3]), .Y(n354) );
  OAI21X1 U615 ( .A(n6604), .B(n6875), .C(n358), .Y(n2798) );
  NAND2X1 U616 ( .A(\Mem[16][0] ), .B(n6878), .Y(n358) );
  OAI21X1 U617 ( .A(n6549), .B(n6874), .C(n359), .Y(n2799) );
  NAND2X1 U618 ( .A(\Mem[16][1] ), .B(n6878), .Y(n359) );
  OAI21X1 U619 ( .A(n6494), .B(n6874), .C(n360), .Y(n2800) );
  NAND2X1 U620 ( .A(\Mem[16][2] ), .B(n6878), .Y(n360) );
  OAI21X1 U621 ( .A(n6479), .B(n6874), .C(n361), .Y(n2801) );
  NAND2X1 U622 ( .A(\Mem[16][3] ), .B(n6877), .Y(n361) );
  OAI21X1 U623 ( .A(n6474), .B(n6874), .C(n362), .Y(n2802) );
  NAND2X1 U624 ( .A(\Mem[16][4] ), .B(n6878), .Y(n362) );
  OAI21X1 U625 ( .A(n6469), .B(n6874), .C(n363), .Y(n2803) );
  NAND2X1 U626 ( .A(\Mem[16][5] ), .B(n6877), .Y(n363) );
  OAI21X1 U627 ( .A(n6464), .B(n6874), .C(n364), .Y(n2804) );
  NAND2X1 U628 ( .A(\Mem[16][6] ), .B(n6877), .Y(n364) );
  OAI21X1 U629 ( .A(n6459), .B(n6874), .C(n365), .Y(n2805) );
  NAND2X1 U630 ( .A(\Mem[16][7] ), .B(n6877), .Y(n365) );
  OAI21X1 U631 ( .A(n6454), .B(n6874), .C(n366), .Y(n2806) );
  NAND2X1 U632 ( .A(\Mem[16][8] ), .B(n6877), .Y(n366) );
  OAI21X1 U633 ( .A(n6449), .B(n6874), .C(n367), .Y(n2807) );
  NAND2X1 U634 ( .A(\Mem[16][9] ), .B(n6877), .Y(n367) );
  OAI21X1 U635 ( .A(n6599), .B(n6874), .C(n368), .Y(n2808) );
  NAND2X1 U636 ( .A(\Mem[16][10] ), .B(n6877), .Y(n368) );
  OAI21X1 U637 ( .A(n6594), .B(n6874), .C(n369), .Y(n2809) );
  NAND2X1 U638 ( .A(\Mem[16][11] ), .B(n6877), .Y(n369) );
  OAI21X1 U639 ( .A(n6589), .B(n6874), .C(n370), .Y(n2810) );
  NAND2X1 U640 ( .A(\Mem[16][12] ), .B(n6877), .Y(n370) );
  OAI21X1 U641 ( .A(n6584), .B(n6875), .C(n371), .Y(n2811) );
  NAND2X1 U642 ( .A(\Mem[16][13] ), .B(n6877), .Y(n371) );
  OAI21X1 U643 ( .A(n6579), .B(n6875), .C(n372), .Y(n2812) );
  NAND2X1 U644 ( .A(\Mem[16][14] ), .B(n6877), .Y(n372) );
  OAI21X1 U645 ( .A(n6574), .B(n6875), .C(n373), .Y(n2813) );
  NAND2X1 U646 ( .A(\Mem[16][15] ), .B(n6876), .Y(n373) );
  OAI21X1 U647 ( .A(n6569), .B(n6875), .C(n374), .Y(n2814) );
  NAND2X1 U648 ( .A(\Mem[16][16] ), .B(n6877), .Y(n374) );
  OAI21X1 U649 ( .A(n6564), .B(n6875), .C(n375), .Y(n2815) );
  NAND2X1 U650 ( .A(\Mem[16][17] ), .B(n6876), .Y(n375) );
  OAI21X1 U651 ( .A(n6559), .B(n6875), .C(n376), .Y(n2816) );
  NAND2X1 U652 ( .A(\Mem[16][18] ), .B(n6876), .Y(n376) );
  OAI21X1 U653 ( .A(n6554), .B(n6875), .C(n377), .Y(n2817) );
  NAND2X1 U654 ( .A(\Mem[16][19] ), .B(n6876), .Y(n377) );
  OAI21X1 U655 ( .A(n6544), .B(n6875), .C(n378), .Y(n2818) );
  NAND2X1 U656 ( .A(\Mem[16][20] ), .B(n6876), .Y(n378) );
  OAI21X1 U657 ( .A(n6539), .B(n6875), .C(n379), .Y(n2819) );
  NAND2X1 U658 ( .A(\Mem[16][21] ), .B(n6876), .Y(n379) );
  OAI21X1 U659 ( .A(n6534), .B(n6875), .C(n380), .Y(n2820) );
  NAND2X1 U660 ( .A(\Mem[16][22] ), .B(n6877), .Y(n380) );
  OAI21X1 U661 ( .A(n6529), .B(n6876), .C(n381), .Y(n2821) );
  NAND2X1 U662 ( .A(\Mem[16][23] ), .B(n6876), .Y(n381) );
  OAI21X1 U663 ( .A(n6524), .B(n6875), .C(n382), .Y(n2822) );
  NAND2X1 U664 ( .A(\Mem[16][24] ), .B(n6877), .Y(n382) );
  OAI21X1 U665 ( .A(n6519), .B(n6876), .C(n383), .Y(n2823) );
  NAND2X1 U666 ( .A(\Mem[16][25] ), .B(n6877), .Y(n383) );
  OAI21X1 U667 ( .A(n6514), .B(n6876), .C(n384), .Y(n2824) );
  NAND2X1 U668 ( .A(\Mem[16][26] ), .B(n6877), .Y(n384) );
  OAI21X1 U669 ( .A(n6509), .B(n6876), .C(n385), .Y(n2825) );
  NAND2X1 U670 ( .A(\Mem[16][27] ), .B(n6877), .Y(n385) );
  OAI21X1 U671 ( .A(n6504), .B(n6876), .C(n386), .Y(n2826) );
  NAND2X1 U672 ( .A(\Mem[16][28] ), .B(n6877), .Y(n386) );
  OAI21X1 U673 ( .A(n6499), .B(n6876), .C(n387), .Y(n2827) );
  NAND2X1 U674 ( .A(\Mem[16][29] ), .B(n6877), .Y(n387) );
  OAI21X1 U675 ( .A(n6489), .B(n6876), .C(n388), .Y(n2828) );
  NAND2X1 U676 ( .A(\Mem[16][30] ), .B(n6878), .Y(n388) );
  OAI21X1 U677 ( .A(n6484), .B(n6876), .C(n389), .Y(n2829) );
  NAND2X1 U678 ( .A(\Mem[16][31] ), .B(n6878), .Y(n389) );
  NAND2X1 U679 ( .A(n7006), .B(n7016), .Y(n357) );
  OAI21X1 U680 ( .A(n6604), .B(n6870), .C(n392), .Y(n2830) );
  NAND2X1 U681 ( .A(\Mem[17][0] ), .B(n6873), .Y(n392) );
  OAI21X1 U682 ( .A(n6549), .B(n6869), .C(n393), .Y(n2831) );
  NAND2X1 U683 ( .A(\Mem[17][1] ), .B(n6873), .Y(n393) );
  OAI21X1 U684 ( .A(n6494), .B(n6869), .C(n394), .Y(n2832) );
  NAND2X1 U685 ( .A(\Mem[17][2] ), .B(n6873), .Y(n394) );
  OAI21X1 U686 ( .A(n6479), .B(n6869), .C(n395), .Y(n2833) );
  NAND2X1 U687 ( .A(\Mem[17][3] ), .B(n6872), .Y(n395) );
  OAI21X1 U688 ( .A(n6474), .B(n6869), .C(n396), .Y(n2834) );
  NAND2X1 U689 ( .A(\Mem[17][4] ), .B(n6873), .Y(n396) );
  OAI21X1 U690 ( .A(n6469), .B(n6869), .C(n397), .Y(n2835) );
  NAND2X1 U691 ( .A(\Mem[17][5] ), .B(n6872), .Y(n397) );
  OAI21X1 U692 ( .A(n6464), .B(n6869), .C(n398), .Y(n2836) );
  NAND2X1 U693 ( .A(\Mem[17][6] ), .B(n6872), .Y(n398) );
  OAI21X1 U694 ( .A(n6459), .B(n6869), .C(n399), .Y(n2837) );
  NAND2X1 U695 ( .A(\Mem[17][7] ), .B(n6872), .Y(n399) );
  OAI21X1 U696 ( .A(n6454), .B(n6869), .C(n400), .Y(n2838) );
  NAND2X1 U697 ( .A(\Mem[17][8] ), .B(n6872), .Y(n400) );
  OAI21X1 U698 ( .A(n6449), .B(n6869), .C(n401), .Y(n2839) );
  NAND2X1 U699 ( .A(\Mem[17][9] ), .B(n6872), .Y(n401) );
  OAI21X1 U700 ( .A(n6599), .B(n6869), .C(n402), .Y(n2840) );
  NAND2X1 U701 ( .A(\Mem[17][10] ), .B(n6872), .Y(n402) );
  OAI21X1 U702 ( .A(n6594), .B(n6869), .C(n403), .Y(n2841) );
  NAND2X1 U703 ( .A(\Mem[17][11] ), .B(n6872), .Y(n403) );
  OAI21X1 U704 ( .A(n6589), .B(n6869), .C(n404), .Y(n2842) );
  NAND2X1 U705 ( .A(\Mem[17][12] ), .B(n6872), .Y(n404) );
  OAI21X1 U706 ( .A(n6584), .B(n6870), .C(n405), .Y(n2843) );
  NAND2X1 U707 ( .A(\Mem[17][13] ), .B(n6872), .Y(n405) );
  OAI21X1 U708 ( .A(n6579), .B(n6870), .C(n406), .Y(n2844) );
  NAND2X1 U709 ( .A(\Mem[17][14] ), .B(n6872), .Y(n406) );
  OAI21X1 U710 ( .A(n6574), .B(n6870), .C(n407), .Y(n2845) );
  NAND2X1 U711 ( .A(\Mem[17][15] ), .B(n6871), .Y(n407) );
  OAI21X1 U712 ( .A(n6569), .B(n6870), .C(n408), .Y(n2846) );
  NAND2X1 U713 ( .A(\Mem[17][16] ), .B(n6872), .Y(n408) );
  OAI21X1 U714 ( .A(n6564), .B(n6870), .C(n409), .Y(n2847) );
  NAND2X1 U715 ( .A(\Mem[17][17] ), .B(n6871), .Y(n409) );
  OAI21X1 U716 ( .A(n6559), .B(n6870), .C(n410), .Y(n2848) );
  NAND2X1 U717 ( .A(\Mem[17][18] ), .B(n6871), .Y(n410) );
  OAI21X1 U718 ( .A(n6554), .B(n6870), .C(n411), .Y(n2849) );
  NAND2X1 U719 ( .A(\Mem[17][19] ), .B(n6871), .Y(n411) );
  OAI21X1 U720 ( .A(n6544), .B(n6870), .C(n412), .Y(n2850) );
  NAND2X1 U721 ( .A(\Mem[17][20] ), .B(n6871), .Y(n412) );
  OAI21X1 U722 ( .A(n6539), .B(n6870), .C(n413), .Y(n2851) );
  NAND2X1 U723 ( .A(\Mem[17][21] ), .B(n6871), .Y(n413) );
  OAI21X1 U724 ( .A(n6534), .B(n6870), .C(n414), .Y(n2852) );
  NAND2X1 U725 ( .A(\Mem[17][22] ), .B(n6872), .Y(n414) );
  OAI21X1 U726 ( .A(n6529), .B(n6871), .C(n415), .Y(n2853) );
  NAND2X1 U727 ( .A(\Mem[17][23] ), .B(n6871), .Y(n415) );
  OAI21X1 U728 ( .A(n6524), .B(n6870), .C(n416), .Y(n2854) );
  NAND2X1 U729 ( .A(\Mem[17][24] ), .B(n6872), .Y(n416) );
  OAI21X1 U730 ( .A(n6519), .B(n6871), .C(n417), .Y(n2855) );
  NAND2X1 U731 ( .A(\Mem[17][25] ), .B(n6872), .Y(n417) );
  OAI21X1 U732 ( .A(n6514), .B(n6871), .C(n418), .Y(n2856) );
  NAND2X1 U733 ( .A(\Mem[17][26] ), .B(n6872), .Y(n418) );
  OAI21X1 U734 ( .A(n6509), .B(n6871), .C(n419), .Y(n2857) );
  NAND2X1 U735 ( .A(\Mem[17][27] ), .B(n6872), .Y(n419) );
  OAI21X1 U736 ( .A(n6504), .B(n6871), .C(n420), .Y(n2858) );
  NAND2X1 U737 ( .A(\Mem[17][28] ), .B(n6872), .Y(n420) );
  OAI21X1 U738 ( .A(n6499), .B(n6871), .C(n421), .Y(n2859) );
  NAND2X1 U739 ( .A(\Mem[17][29] ), .B(n6872), .Y(n421) );
  OAI21X1 U740 ( .A(n6489), .B(n6871), .C(n422), .Y(n2860) );
  NAND2X1 U741 ( .A(\Mem[17][30] ), .B(n6873), .Y(n422) );
  OAI21X1 U742 ( .A(n6484), .B(n6871), .C(n423), .Y(n2861) );
  NAND2X1 U743 ( .A(\Mem[17][31] ), .B(n6873), .Y(n423) );
  NAND2X1 U744 ( .A(n7006), .B(n7017), .Y(n391) );
  OAI21X1 U745 ( .A(n6604), .B(n6865), .C(n425), .Y(n2862) );
  NAND2X1 U746 ( .A(\Mem[18][0] ), .B(n6868), .Y(n425) );
  OAI21X1 U747 ( .A(n6549), .B(n6864), .C(n426), .Y(n2863) );
  NAND2X1 U748 ( .A(\Mem[18][1] ), .B(n6868), .Y(n426) );
  OAI21X1 U749 ( .A(n6494), .B(n6864), .C(n427), .Y(n2864) );
  NAND2X1 U750 ( .A(\Mem[18][2] ), .B(n6868), .Y(n427) );
  OAI21X1 U751 ( .A(n6479), .B(n6864), .C(n428), .Y(n2865) );
  NAND2X1 U752 ( .A(\Mem[18][3] ), .B(n6867), .Y(n428) );
  OAI21X1 U753 ( .A(n6474), .B(n6864), .C(n429), .Y(n2866) );
  NAND2X1 U754 ( .A(\Mem[18][4] ), .B(n6868), .Y(n429) );
  OAI21X1 U755 ( .A(n6469), .B(n6864), .C(n430), .Y(n2867) );
  NAND2X1 U756 ( .A(\Mem[18][5] ), .B(n6867), .Y(n430) );
  OAI21X1 U757 ( .A(n6464), .B(n6864), .C(n431), .Y(n2868) );
  NAND2X1 U758 ( .A(\Mem[18][6] ), .B(n6867), .Y(n431) );
  OAI21X1 U759 ( .A(n6459), .B(n6864), .C(n432), .Y(n2869) );
  NAND2X1 U760 ( .A(\Mem[18][7] ), .B(n6867), .Y(n432) );
  OAI21X1 U761 ( .A(n6454), .B(n6864), .C(n433), .Y(n2870) );
  NAND2X1 U762 ( .A(\Mem[18][8] ), .B(n6867), .Y(n433) );
  OAI21X1 U763 ( .A(n6449), .B(n6864), .C(n434), .Y(n2871) );
  NAND2X1 U764 ( .A(\Mem[18][9] ), .B(n6867), .Y(n434) );
  OAI21X1 U765 ( .A(n6599), .B(n6864), .C(n435), .Y(n2872) );
  NAND2X1 U766 ( .A(\Mem[18][10] ), .B(n6867), .Y(n435) );
  OAI21X1 U767 ( .A(n6594), .B(n6864), .C(n436), .Y(n2873) );
  NAND2X1 U768 ( .A(\Mem[18][11] ), .B(n6867), .Y(n436) );
  OAI21X1 U769 ( .A(n6589), .B(n6864), .C(n437), .Y(n2874) );
  NAND2X1 U770 ( .A(\Mem[18][12] ), .B(n6867), .Y(n437) );
  OAI21X1 U771 ( .A(n6584), .B(n6865), .C(n438), .Y(n2875) );
  NAND2X1 U772 ( .A(\Mem[18][13] ), .B(n6867), .Y(n438) );
  OAI21X1 U773 ( .A(n6579), .B(n6865), .C(n439), .Y(n2876) );
  NAND2X1 U774 ( .A(\Mem[18][14] ), .B(n6867), .Y(n439) );
  OAI21X1 U775 ( .A(n6574), .B(n6865), .C(n440), .Y(n2877) );
  NAND2X1 U776 ( .A(\Mem[18][15] ), .B(n6866), .Y(n440) );
  OAI21X1 U777 ( .A(n6569), .B(n6865), .C(n441), .Y(n2878) );
  NAND2X1 U778 ( .A(\Mem[18][16] ), .B(n6867), .Y(n441) );
  OAI21X1 U779 ( .A(n6564), .B(n6865), .C(n442), .Y(n2879) );
  NAND2X1 U780 ( .A(\Mem[18][17] ), .B(n6866), .Y(n442) );
  OAI21X1 U781 ( .A(n6559), .B(n6865), .C(n443), .Y(n2880) );
  NAND2X1 U782 ( .A(\Mem[18][18] ), .B(n6866), .Y(n443) );
  OAI21X1 U783 ( .A(n6554), .B(n6865), .C(n444), .Y(n2881) );
  NAND2X1 U784 ( .A(\Mem[18][19] ), .B(n6866), .Y(n444) );
  OAI21X1 U785 ( .A(n6544), .B(n6865), .C(n445), .Y(n2882) );
  NAND2X1 U786 ( .A(\Mem[18][20] ), .B(n6866), .Y(n445) );
  OAI21X1 U787 ( .A(n6539), .B(n6865), .C(n446), .Y(n2883) );
  NAND2X1 U788 ( .A(\Mem[18][21] ), .B(n6866), .Y(n446) );
  OAI21X1 U789 ( .A(n6534), .B(n6865), .C(n447), .Y(n2884) );
  NAND2X1 U790 ( .A(\Mem[18][22] ), .B(n6867), .Y(n447) );
  OAI21X1 U791 ( .A(n6529), .B(n6866), .C(n448), .Y(n2885) );
  NAND2X1 U792 ( .A(\Mem[18][23] ), .B(n6866), .Y(n448) );
  OAI21X1 U793 ( .A(n6524), .B(n6865), .C(n449), .Y(n2886) );
  NAND2X1 U794 ( .A(\Mem[18][24] ), .B(n6867), .Y(n449) );
  OAI21X1 U795 ( .A(n6519), .B(n6866), .C(n450), .Y(n2887) );
  NAND2X1 U796 ( .A(\Mem[18][25] ), .B(n6867), .Y(n450) );
  OAI21X1 U797 ( .A(n6514), .B(n6866), .C(n451), .Y(n2888) );
  NAND2X1 U798 ( .A(\Mem[18][26] ), .B(n6867), .Y(n451) );
  OAI21X1 U799 ( .A(n6509), .B(n6866), .C(n452), .Y(n2889) );
  NAND2X1 U800 ( .A(\Mem[18][27] ), .B(n6867), .Y(n452) );
  OAI21X1 U801 ( .A(n6504), .B(n6866), .C(n453), .Y(n2890) );
  NAND2X1 U802 ( .A(\Mem[18][28] ), .B(n6867), .Y(n453) );
  OAI21X1 U803 ( .A(n6499), .B(n6866), .C(n454), .Y(n2891) );
  NAND2X1 U804 ( .A(\Mem[18][29] ), .B(n6867), .Y(n454) );
  OAI21X1 U805 ( .A(n6489), .B(n6866), .C(n455), .Y(n2892) );
  NAND2X1 U806 ( .A(\Mem[18][30] ), .B(n6868), .Y(n455) );
  OAI21X1 U807 ( .A(n6484), .B(n6866), .C(n456), .Y(n2893) );
  NAND2X1 U808 ( .A(\Mem[18][31] ), .B(n6868), .Y(n456) );
  NAND2X1 U809 ( .A(n7006), .B(n7018), .Y(n424) );
  OAI21X1 U810 ( .A(n6605), .B(n6860), .C(n458), .Y(n2894) );
  NAND2X1 U811 ( .A(\Mem[19][0] ), .B(n6863), .Y(n458) );
  OAI21X1 U812 ( .A(n6550), .B(n6859), .C(n459), .Y(n2895) );
  NAND2X1 U813 ( .A(\Mem[19][1] ), .B(n6863), .Y(n459) );
  OAI21X1 U814 ( .A(n6495), .B(n6859), .C(n460), .Y(n2896) );
  NAND2X1 U815 ( .A(\Mem[19][2] ), .B(n6863), .Y(n460) );
  OAI21X1 U816 ( .A(n6480), .B(n6859), .C(n461), .Y(n2897) );
  NAND2X1 U817 ( .A(\Mem[19][3] ), .B(n6862), .Y(n461) );
  OAI21X1 U818 ( .A(n6475), .B(n6859), .C(n462), .Y(n2898) );
  NAND2X1 U819 ( .A(\Mem[19][4] ), .B(n6863), .Y(n462) );
  OAI21X1 U820 ( .A(n6470), .B(n6859), .C(n463), .Y(n2899) );
  NAND2X1 U821 ( .A(\Mem[19][5] ), .B(n6862), .Y(n463) );
  OAI21X1 U822 ( .A(n6465), .B(n6859), .C(n464), .Y(n2900) );
  NAND2X1 U823 ( .A(\Mem[19][6] ), .B(n6862), .Y(n464) );
  OAI21X1 U824 ( .A(n6460), .B(n6859), .C(n465), .Y(n2901) );
  NAND2X1 U825 ( .A(\Mem[19][7] ), .B(n6862), .Y(n465) );
  OAI21X1 U826 ( .A(n6455), .B(n6859), .C(n466), .Y(n2902) );
  NAND2X1 U827 ( .A(\Mem[19][8] ), .B(n6862), .Y(n466) );
  OAI21X1 U828 ( .A(n6450), .B(n6859), .C(n467), .Y(n2903) );
  NAND2X1 U829 ( .A(\Mem[19][9] ), .B(n6862), .Y(n467) );
  OAI21X1 U830 ( .A(n6600), .B(n6859), .C(n468), .Y(n2904) );
  NAND2X1 U831 ( .A(\Mem[19][10] ), .B(n6862), .Y(n468) );
  OAI21X1 U832 ( .A(n6595), .B(n6859), .C(n469), .Y(n2905) );
  NAND2X1 U833 ( .A(\Mem[19][11] ), .B(n6862), .Y(n469) );
  OAI21X1 U834 ( .A(n6590), .B(n6859), .C(n470), .Y(n2906) );
  NAND2X1 U835 ( .A(\Mem[19][12] ), .B(n6862), .Y(n470) );
  OAI21X1 U836 ( .A(n6585), .B(n6860), .C(n471), .Y(n2907) );
  NAND2X1 U837 ( .A(\Mem[19][13] ), .B(n6862), .Y(n471) );
  OAI21X1 U838 ( .A(n6580), .B(n6860), .C(n472), .Y(n2908) );
  NAND2X1 U839 ( .A(\Mem[19][14] ), .B(n6862), .Y(n472) );
  OAI21X1 U840 ( .A(n6575), .B(n6860), .C(n473), .Y(n2909) );
  NAND2X1 U841 ( .A(\Mem[19][15] ), .B(n6861), .Y(n473) );
  OAI21X1 U842 ( .A(n6570), .B(n6860), .C(n474), .Y(n2910) );
  NAND2X1 U843 ( .A(\Mem[19][16] ), .B(n6862), .Y(n474) );
  OAI21X1 U844 ( .A(n6565), .B(n6860), .C(n475), .Y(n2911) );
  NAND2X1 U845 ( .A(\Mem[19][17] ), .B(n6861), .Y(n475) );
  OAI21X1 U846 ( .A(n6560), .B(n6860), .C(n476), .Y(n2912) );
  NAND2X1 U847 ( .A(\Mem[19][18] ), .B(n6861), .Y(n476) );
  OAI21X1 U848 ( .A(n6555), .B(n6860), .C(n477), .Y(n2913) );
  NAND2X1 U849 ( .A(\Mem[19][19] ), .B(n6861), .Y(n477) );
  OAI21X1 U850 ( .A(n6545), .B(n6860), .C(n478), .Y(n2914) );
  NAND2X1 U851 ( .A(\Mem[19][20] ), .B(n6861), .Y(n478) );
  OAI21X1 U852 ( .A(n6540), .B(n6860), .C(n479), .Y(n2915) );
  NAND2X1 U853 ( .A(\Mem[19][21] ), .B(n6861), .Y(n479) );
  OAI21X1 U854 ( .A(n6535), .B(n6860), .C(n480), .Y(n2916) );
  NAND2X1 U855 ( .A(\Mem[19][22] ), .B(n6862), .Y(n480) );
  OAI21X1 U856 ( .A(n6530), .B(n6861), .C(n481), .Y(n2917) );
  NAND2X1 U857 ( .A(\Mem[19][23] ), .B(n6861), .Y(n481) );
  OAI21X1 U858 ( .A(n6525), .B(n6860), .C(n482), .Y(n2918) );
  NAND2X1 U859 ( .A(\Mem[19][24] ), .B(n6862), .Y(n482) );
  OAI21X1 U860 ( .A(n6520), .B(n6861), .C(n483), .Y(n2919) );
  NAND2X1 U861 ( .A(\Mem[19][25] ), .B(n6862), .Y(n483) );
  OAI21X1 U862 ( .A(n6515), .B(n6861), .C(n484), .Y(n2920) );
  NAND2X1 U863 ( .A(\Mem[19][26] ), .B(n6862), .Y(n484) );
  OAI21X1 U864 ( .A(n6510), .B(n6861), .C(n485), .Y(n2921) );
  NAND2X1 U865 ( .A(\Mem[19][27] ), .B(n6862), .Y(n485) );
  OAI21X1 U866 ( .A(n6505), .B(n6861), .C(n486), .Y(n2922) );
  NAND2X1 U867 ( .A(\Mem[19][28] ), .B(n6862), .Y(n486) );
  OAI21X1 U868 ( .A(n6500), .B(n6861), .C(n487), .Y(n2923) );
  NAND2X1 U869 ( .A(\Mem[19][29] ), .B(n6862), .Y(n487) );
  OAI21X1 U870 ( .A(n6490), .B(n6861), .C(n488), .Y(n2924) );
  NAND2X1 U871 ( .A(\Mem[19][30] ), .B(n6863), .Y(n488) );
  OAI21X1 U872 ( .A(n6485), .B(n6861), .C(n489), .Y(n2925) );
  NAND2X1 U873 ( .A(\Mem[19][31] ), .B(n6863), .Y(n489) );
  NAND2X1 U874 ( .A(n7006), .B(n7019), .Y(n457) );
  OAI21X1 U875 ( .A(n6605), .B(n6855), .C(n491), .Y(n2926) );
  NAND2X1 U876 ( .A(\Mem[20][0] ), .B(n6858), .Y(n491) );
  OAI21X1 U877 ( .A(n6550), .B(n6854), .C(n492), .Y(n2927) );
  NAND2X1 U878 ( .A(\Mem[20][1] ), .B(n6858), .Y(n492) );
  OAI21X1 U879 ( .A(n6495), .B(n6854), .C(n493), .Y(n2928) );
  NAND2X1 U880 ( .A(\Mem[20][2] ), .B(n6858), .Y(n493) );
  OAI21X1 U881 ( .A(n6480), .B(n6854), .C(n494), .Y(n2929) );
  NAND2X1 U882 ( .A(\Mem[20][3] ), .B(n6857), .Y(n494) );
  OAI21X1 U883 ( .A(n6475), .B(n6854), .C(n495), .Y(n2930) );
  NAND2X1 U884 ( .A(\Mem[20][4] ), .B(n6858), .Y(n495) );
  OAI21X1 U885 ( .A(n6470), .B(n6854), .C(n496), .Y(n2931) );
  NAND2X1 U886 ( .A(\Mem[20][5] ), .B(n6857), .Y(n496) );
  OAI21X1 U887 ( .A(n6465), .B(n6854), .C(n497), .Y(n2932) );
  NAND2X1 U888 ( .A(\Mem[20][6] ), .B(n6857), .Y(n497) );
  OAI21X1 U889 ( .A(n6460), .B(n6854), .C(n498), .Y(n2933) );
  NAND2X1 U890 ( .A(\Mem[20][7] ), .B(n6857), .Y(n498) );
  OAI21X1 U891 ( .A(n6455), .B(n6854), .C(n499), .Y(n2934) );
  NAND2X1 U892 ( .A(\Mem[20][8] ), .B(n6857), .Y(n499) );
  OAI21X1 U893 ( .A(n6450), .B(n6854), .C(n500), .Y(n2935) );
  NAND2X1 U894 ( .A(\Mem[20][9] ), .B(n6857), .Y(n500) );
  OAI21X1 U895 ( .A(n6600), .B(n6854), .C(n501), .Y(n2936) );
  NAND2X1 U896 ( .A(\Mem[20][10] ), .B(n6857), .Y(n501) );
  OAI21X1 U897 ( .A(n6595), .B(n6854), .C(n502), .Y(n2937) );
  NAND2X1 U898 ( .A(\Mem[20][11] ), .B(n6857), .Y(n502) );
  OAI21X1 U899 ( .A(n6590), .B(n6854), .C(n503), .Y(n2938) );
  NAND2X1 U900 ( .A(\Mem[20][12] ), .B(n6857), .Y(n503) );
  OAI21X1 U901 ( .A(n6585), .B(n6855), .C(n504), .Y(n2939) );
  NAND2X1 U902 ( .A(\Mem[20][13] ), .B(n6857), .Y(n504) );
  OAI21X1 U903 ( .A(n6580), .B(n6855), .C(n505), .Y(n2940) );
  NAND2X1 U904 ( .A(\Mem[20][14] ), .B(n6857), .Y(n505) );
  OAI21X1 U905 ( .A(n6575), .B(n6855), .C(n506), .Y(n2941) );
  NAND2X1 U906 ( .A(\Mem[20][15] ), .B(n6856), .Y(n506) );
  OAI21X1 U907 ( .A(n6570), .B(n6855), .C(n507), .Y(n2942) );
  NAND2X1 U908 ( .A(\Mem[20][16] ), .B(n6857), .Y(n507) );
  OAI21X1 U909 ( .A(n6565), .B(n6855), .C(n508), .Y(n2943) );
  NAND2X1 U910 ( .A(\Mem[20][17] ), .B(n6856), .Y(n508) );
  OAI21X1 U911 ( .A(n6560), .B(n6855), .C(n509), .Y(n2944) );
  NAND2X1 U912 ( .A(\Mem[20][18] ), .B(n6856), .Y(n509) );
  OAI21X1 U913 ( .A(n6555), .B(n6855), .C(n510), .Y(n2945) );
  NAND2X1 U914 ( .A(\Mem[20][19] ), .B(n6856), .Y(n510) );
  OAI21X1 U915 ( .A(n6545), .B(n6855), .C(n511), .Y(n2946) );
  NAND2X1 U916 ( .A(\Mem[20][20] ), .B(n6856), .Y(n511) );
  OAI21X1 U917 ( .A(n6540), .B(n6855), .C(n512), .Y(n2947) );
  NAND2X1 U918 ( .A(\Mem[20][21] ), .B(n6856), .Y(n512) );
  OAI21X1 U919 ( .A(n6535), .B(n6855), .C(n513), .Y(n2948) );
  NAND2X1 U920 ( .A(\Mem[20][22] ), .B(n6857), .Y(n513) );
  OAI21X1 U921 ( .A(n6530), .B(n6856), .C(n514), .Y(n2949) );
  NAND2X1 U922 ( .A(\Mem[20][23] ), .B(n6856), .Y(n514) );
  OAI21X1 U923 ( .A(n6525), .B(n6855), .C(n515), .Y(n2950) );
  NAND2X1 U924 ( .A(\Mem[20][24] ), .B(n6857), .Y(n515) );
  OAI21X1 U925 ( .A(n6520), .B(n6856), .C(n516), .Y(n2951) );
  NAND2X1 U926 ( .A(\Mem[20][25] ), .B(n6857), .Y(n516) );
  OAI21X1 U927 ( .A(n6515), .B(n6856), .C(n517), .Y(n2952) );
  NAND2X1 U928 ( .A(\Mem[20][26] ), .B(n6857), .Y(n517) );
  OAI21X1 U929 ( .A(n6510), .B(n6856), .C(n518), .Y(n2953) );
  NAND2X1 U930 ( .A(\Mem[20][27] ), .B(n6857), .Y(n518) );
  OAI21X1 U931 ( .A(n6505), .B(n6856), .C(n519), .Y(n2954) );
  NAND2X1 U932 ( .A(\Mem[20][28] ), .B(n6857), .Y(n519) );
  OAI21X1 U933 ( .A(n6500), .B(n6856), .C(n520), .Y(n2955) );
  NAND2X1 U934 ( .A(\Mem[20][29] ), .B(n6857), .Y(n520) );
  OAI21X1 U935 ( .A(n6490), .B(n6856), .C(n521), .Y(n2956) );
  NAND2X1 U936 ( .A(\Mem[20][30] ), .B(n6858), .Y(n521) );
  OAI21X1 U937 ( .A(n6485), .B(n6856), .C(n522), .Y(n2957) );
  NAND2X1 U938 ( .A(\Mem[20][31] ), .B(n6858), .Y(n522) );
  NAND2X1 U939 ( .A(n7006), .B(n7022), .Y(n490) );
  OAI21X1 U940 ( .A(n6605), .B(n6850), .C(n524), .Y(n2958) );
  NAND2X1 U941 ( .A(\Mem[21][0] ), .B(n6853), .Y(n524) );
  OAI21X1 U942 ( .A(n6550), .B(n6849), .C(n525), .Y(n2959) );
  NAND2X1 U943 ( .A(\Mem[21][1] ), .B(n6853), .Y(n525) );
  OAI21X1 U944 ( .A(n6495), .B(n6849), .C(n526), .Y(n2960) );
  NAND2X1 U945 ( .A(\Mem[21][2] ), .B(n6853), .Y(n526) );
  OAI21X1 U946 ( .A(n6480), .B(n6849), .C(n527), .Y(n2961) );
  NAND2X1 U947 ( .A(\Mem[21][3] ), .B(n6852), .Y(n527) );
  OAI21X1 U948 ( .A(n6475), .B(n6849), .C(n528), .Y(n2962) );
  NAND2X1 U949 ( .A(\Mem[21][4] ), .B(n6853), .Y(n528) );
  OAI21X1 U950 ( .A(n6470), .B(n6849), .C(n529), .Y(n2963) );
  NAND2X1 U951 ( .A(\Mem[21][5] ), .B(n6852), .Y(n529) );
  OAI21X1 U952 ( .A(n6465), .B(n6849), .C(n530), .Y(n2964) );
  NAND2X1 U953 ( .A(\Mem[21][6] ), .B(n6852), .Y(n530) );
  OAI21X1 U954 ( .A(n6460), .B(n6849), .C(n531), .Y(n2965) );
  NAND2X1 U955 ( .A(\Mem[21][7] ), .B(n6852), .Y(n531) );
  OAI21X1 U956 ( .A(n6455), .B(n6849), .C(n532), .Y(n2966) );
  NAND2X1 U957 ( .A(\Mem[21][8] ), .B(n6852), .Y(n532) );
  OAI21X1 U958 ( .A(n6450), .B(n6849), .C(n533), .Y(n2967) );
  NAND2X1 U959 ( .A(\Mem[21][9] ), .B(n6852), .Y(n533) );
  OAI21X1 U960 ( .A(n6600), .B(n6849), .C(n534), .Y(n2968) );
  NAND2X1 U961 ( .A(\Mem[21][10] ), .B(n6852), .Y(n534) );
  OAI21X1 U962 ( .A(n6595), .B(n6849), .C(n535), .Y(n2969) );
  NAND2X1 U963 ( .A(\Mem[21][11] ), .B(n6852), .Y(n535) );
  OAI21X1 U964 ( .A(n6590), .B(n6849), .C(n536), .Y(n2970) );
  NAND2X1 U965 ( .A(\Mem[21][12] ), .B(n6852), .Y(n536) );
  OAI21X1 U966 ( .A(n6585), .B(n6850), .C(n537), .Y(n2971) );
  NAND2X1 U967 ( .A(\Mem[21][13] ), .B(n6852), .Y(n537) );
  OAI21X1 U968 ( .A(n6580), .B(n6850), .C(n538), .Y(n2972) );
  NAND2X1 U969 ( .A(\Mem[21][14] ), .B(n6852), .Y(n538) );
  OAI21X1 U970 ( .A(n6575), .B(n6850), .C(n539), .Y(n2973) );
  NAND2X1 U971 ( .A(\Mem[21][15] ), .B(n6851), .Y(n539) );
  OAI21X1 U972 ( .A(n6570), .B(n6850), .C(n540), .Y(n2974) );
  NAND2X1 U973 ( .A(\Mem[21][16] ), .B(n6852), .Y(n540) );
  OAI21X1 U974 ( .A(n6565), .B(n6850), .C(n541), .Y(n2975) );
  NAND2X1 U975 ( .A(\Mem[21][17] ), .B(n6851), .Y(n541) );
  OAI21X1 U976 ( .A(n6560), .B(n6850), .C(n542), .Y(n2976) );
  NAND2X1 U977 ( .A(\Mem[21][18] ), .B(n6851), .Y(n542) );
  OAI21X1 U978 ( .A(n6555), .B(n6850), .C(n543), .Y(n2977) );
  NAND2X1 U979 ( .A(\Mem[21][19] ), .B(n6851), .Y(n543) );
  OAI21X1 U980 ( .A(n6545), .B(n6850), .C(n544), .Y(n2978) );
  NAND2X1 U981 ( .A(\Mem[21][20] ), .B(n6851), .Y(n544) );
  OAI21X1 U982 ( .A(n6540), .B(n6850), .C(n545), .Y(n2979) );
  NAND2X1 U983 ( .A(\Mem[21][21] ), .B(n6851), .Y(n545) );
  OAI21X1 U984 ( .A(n6535), .B(n6850), .C(n546), .Y(n2980) );
  NAND2X1 U985 ( .A(\Mem[21][22] ), .B(n6852), .Y(n546) );
  OAI21X1 U986 ( .A(n6530), .B(n6851), .C(n547), .Y(n2981) );
  NAND2X1 U987 ( .A(\Mem[21][23] ), .B(n6851), .Y(n547) );
  OAI21X1 U988 ( .A(n6525), .B(n6850), .C(n548), .Y(n2982) );
  NAND2X1 U989 ( .A(\Mem[21][24] ), .B(n6852), .Y(n548) );
  OAI21X1 U990 ( .A(n6520), .B(n6851), .C(n549), .Y(n2983) );
  NAND2X1 U991 ( .A(\Mem[21][25] ), .B(n6852), .Y(n549) );
  OAI21X1 U992 ( .A(n6515), .B(n6851), .C(n550), .Y(n2984) );
  NAND2X1 U993 ( .A(\Mem[21][26] ), .B(n6852), .Y(n550) );
  OAI21X1 U994 ( .A(n6510), .B(n6851), .C(n551), .Y(n2985) );
  NAND2X1 U995 ( .A(\Mem[21][27] ), .B(n6852), .Y(n551) );
  OAI21X1 U996 ( .A(n6505), .B(n6851), .C(n552), .Y(n2986) );
  NAND2X1 U997 ( .A(\Mem[21][28] ), .B(n6852), .Y(n552) );
  OAI21X1 U998 ( .A(n6500), .B(n6851), .C(n553), .Y(n2987) );
  NAND2X1 U999 ( .A(\Mem[21][29] ), .B(n6852), .Y(n553) );
  OAI21X1 U1000 ( .A(n6490), .B(n6851), .C(n554), .Y(n2988) );
  NAND2X1 U1001 ( .A(\Mem[21][30] ), .B(n6853), .Y(n554) );
  OAI21X1 U1002 ( .A(n6485), .B(n6851), .C(n555), .Y(n2989) );
  NAND2X1 U1003 ( .A(\Mem[21][31] ), .B(n6853), .Y(n555) );
  NAND2X1 U1004 ( .A(n7006), .B(n7023), .Y(n523) );
  OAI21X1 U1005 ( .A(n6605), .B(n6845), .C(n557), .Y(n2990) );
  NAND2X1 U1006 ( .A(\Mem[22][0] ), .B(n6848), .Y(n557) );
  OAI21X1 U1007 ( .A(n6550), .B(n6844), .C(n558), .Y(n2991) );
  NAND2X1 U1008 ( .A(\Mem[22][1] ), .B(n6848), .Y(n558) );
  OAI21X1 U1009 ( .A(n6495), .B(n6844), .C(n559), .Y(n2992) );
  NAND2X1 U1010 ( .A(\Mem[22][2] ), .B(n6848), .Y(n559) );
  OAI21X1 U1011 ( .A(n6480), .B(n6844), .C(n560), .Y(n2993) );
  NAND2X1 U1012 ( .A(\Mem[22][3] ), .B(n6847), .Y(n560) );
  OAI21X1 U1013 ( .A(n6475), .B(n6844), .C(n561), .Y(n2994) );
  NAND2X1 U1014 ( .A(\Mem[22][4] ), .B(n6848), .Y(n561) );
  OAI21X1 U1015 ( .A(n6470), .B(n6844), .C(n562), .Y(n2995) );
  NAND2X1 U1016 ( .A(\Mem[22][5] ), .B(n6847), .Y(n562) );
  OAI21X1 U1017 ( .A(n6465), .B(n6844), .C(n563), .Y(n2996) );
  NAND2X1 U1018 ( .A(\Mem[22][6] ), .B(n6847), .Y(n563) );
  OAI21X1 U1019 ( .A(n6460), .B(n6844), .C(n564), .Y(n2997) );
  NAND2X1 U1020 ( .A(\Mem[22][7] ), .B(n6847), .Y(n564) );
  OAI21X1 U1021 ( .A(n6455), .B(n6844), .C(n565), .Y(n2998) );
  NAND2X1 U1022 ( .A(\Mem[22][8] ), .B(n6847), .Y(n565) );
  OAI21X1 U1023 ( .A(n6450), .B(n6844), .C(n566), .Y(n2999) );
  NAND2X1 U1024 ( .A(\Mem[22][9] ), .B(n6847), .Y(n566) );
  OAI21X1 U1025 ( .A(n6600), .B(n6844), .C(n567), .Y(n3000) );
  NAND2X1 U1026 ( .A(\Mem[22][10] ), .B(n6847), .Y(n567) );
  OAI21X1 U1027 ( .A(n6595), .B(n6844), .C(n568), .Y(n3001) );
  NAND2X1 U1028 ( .A(\Mem[22][11] ), .B(n6847), .Y(n568) );
  OAI21X1 U1029 ( .A(n6590), .B(n6844), .C(n569), .Y(n3002) );
  NAND2X1 U1030 ( .A(\Mem[22][12] ), .B(n6847), .Y(n569) );
  OAI21X1 U1031 ( .A(n6585), .B(n6845), .C(n570), .Y(n3003) );
  NAND2X1 U1032 ( .A(\Mem[22][13] ), .B(n6847), .Y(n570) );
  OAI21X1 U1033 ( .A(n6580), .B(n6845), .C(n571), .Y(n3004) );
  NAND2X1 U1034 ( .A(\Mem[22][14] ), .B(n6847), .Y(n571) );
  OAI21X1 U1035 ( .A(n6575), .B(n6845), .C(n572), .Y(n3005) );
  NAND2X1 U1036 ( .A(\Mem[22][15] ), .B(n6846), .Y(n572) );
  OAI21X1 U1037 ( .A(n6570), .B(n6845), .C(n573), .Y(n3006) );
  NAND2X1 U1038 ( .A(\Mem[22][16] ), .B(n6847), .Y(n573) );
  OAI21X1 U1039 ( .A(n6565), .B(n6845), .C(n574), .Y(n3007) );
  NAND2X1 U1040 ( .A(\Mem[22][17] ), .B(n6846), .Y(n574) );
  OAI21X1 U1041 ( .A(n6560), .B(n6845), .C(n575), .Y(n3008) );
  NAND2X1 U1042 ( .A(\Mem[22][18] ), .B(n6846), .Y(n575) );
  OAI21X1 U1043 ( .A(n6555), .B(n6845), .C(n576), .Y(n3009) );
  NAND2X1 U1044 ( .A(\Mem[22][19] ), .B(n6846), .Y(n576) );
  OAI21X1 U1045 ( .A(n6545), .B(n6845), .C(n577), .Y(n3010) );
  NAND2X1 U1046 ( .A(\Mem[22][20] ), .B(n6846), .Y(n577) );
  OAI21X1 U1047 ( .A(n6540), .B(n6845), .C(n578), .Y(n3011) );
  NAND2X1 U1048 ( .A(\Mem[22][21] ), .B(n6846), .Y(n578) );
  OAI21X1 U1049 ( .A(n6535), .B(n6845), .C(n579), .Y(n3012) );
  NAND2X1 U1050 ( .A(\Mem[22][22] ), .B(n6847), .Y(n579) );
  OAI21X1 U1051 ( .A(n6530), .B(n6846), .C(n580), .Y(n3013) );
  NAND2X1 U1052 ( .A(\Mem[22][23] ), .B(n6846), .Y(n580) );
  OAI21X1 U1053 ( .A(n6525), .B(n6845), .C(n581), .Y(n3014) );
  NAND2X1 U1054 ( .A(\Mem[22][24] ), .B(n6847), .Y(n581) );
  OAI21X1 U1055 ( .A(n6520), .B(n6846), .C(n582), .Y(n3015) );
  NAND2X1 U1056 ( .A(\Mem[22][25] ), .B(n6847), .Y(n582) );
  OAI21X1 U1057 ( .A(n6515), .B(n6846), .C(n583), .Y(n3016) );
  NAND2X1 U1058 ( .A(\Mem[22][26] ), .B(n6847), .Y(n583) );
  OAI21X1 U1059 ( .A(n6510), .B(n6846), .C(n584), .Y(n3017) );
  NAND2X1 U1060 ( .A(\Mem[22][27] ), .B(n6847), .Y(n584) );
  OAI21X1 U1061 ( .A(n6505), .B(n6846), .C(n585), .Y(n3018) );
  NAND2X1 U1062 ( .A(\Mem[22][28] ), .B(n6847), .Y(n585) );
  OAI21X1 U1063 ( .A(n6500), .B(n6846), .C(n586), .Y(n3019) );
  NAND2X1 U1064 ( .A(\Mem[22][29] ), .B(n6847), .Y(n586) );
  OAI21X1 U1065 ( .A(n6490), .B(n6846), .C(n587), .Y(n3020) );
  NAND2X1 U1066 ( .A(\Mem[22][30] ), .B(n6848), .Y(n587) );
  OAI21X1 U1067 ( .A(n6485), .B(n6846), .C(n588), .Y(n3021) );
  NAND2X1 U1068 ( .A(\Mem[22][31] ), .B(n6848), .Y(n588) );
  NAND2X1 U1069 ( .A(n7006), .B(n7024), .Y(n556) );
  OAI21X1 U1070 ( .A(n6606), .B(n6840), .C(n590), .Y(n3022) );
  NAND2X1 U1071 ( .A(\Mem[23][0] ), .B(n6843), .Y(n590) );
  OAI21X1 U1072 ( .A(n6551), .B(n6839), .C(n591), .Y(n3023) );
  NAND2X1 U1073 ( .A(\Mem[23][1] ), .B(n6843), .Y(n591) );
  OAI21X1 U1074 ( .A(n6496), .B(n6839), .C(n592), .Y(n3024) );
  NAND2X1 U1075 ( .A(\Mem[23][2] ), .B(n6843), .Y(n592) );
  OAI21X1 U1076 ( .A(n6481), .B(n6839), .C(n593), .Y(n3025) );
  NAND2X1 U1077 ( .A(\Mem[23][3] ), .B(n6842), .Y(n593) );
  OAI21X1 U1078 ( .A(n6476), .B(n6839), .C(n594), .Y(n3026) );
  NAND2X1 U1079 ( .A(\Mem[23][4] ), .B(n6843), .Y(n594) );
  OAI21X1 U1080 ( .A(n6471), .B(n6839), .C(n595), .Y(n3027) );
  NAND2X1 U1081 ( .A(\Mem[23][5] ), .B(n6842), .Y(n595) );
  OAI21X1 U1082 ( .A(n6466), .B(n6839), .C(n596), .Y(n3028) );
  NAND2X1 U1083 ( .A(\Mem[23][6] ), .B(n6842), .Y(n596) );
  OAI21X1 U1084 ( .A(n6461), .B(n6839), .C(n597), .Y(n3029) );
  NAND2X1 U1085 ( .A(\Mem[23][7] ), .B(n6842), .Y(n597) );
  OAI21X1 U1086 ( .A(n6456), .B(n6839), .C(n598), .Y(n3030) );
  NAND2X1 U1087 ( .A(\Mem[23][8] ), .B(n6842), .Y(n598) );
  OAI21X1 U1088 ( .A(n6451), .B(n6839), .C(n599), .Y(n3031) );
  NAND2X1 U1089 ( .A(\Mem[23][9] ), .B(n6842), .Y(n599) );
  OAI21X1 U1090 ( .A(n6601), .B(n6839), .C(n600), .Y(n3032) );
  NAND2X1 U1091 ( .A(\Mem[23][10] ), .B(n6842), .Y(n600) );
  OAI21X1 U1092 ( .A(n6596), .B(n6839), .C(n601), .Y(n3033) );
  NAND2X1 U1093 ( .A(\Mem[23][11] ), .B(n6842), .Y(n601) );
  OAI21X1 U1094 ( .A(n6591), .B(n6839), .C(n602), .Y(n3034) );
  NAND2X1 U1095 ( .A(\Mem[23][12] ), .B(n6842), .Y(n602) );
  OAI21X1 U1096 ( .A(n6586), .B(n6840), .C(n603), .Y(n3035) );
  NAND2X1 U1097 ( .A(\Mem[23][13] ), .B(n6842), .Y(n603) );
  OAI21X1 U1098 ( .A(n6581), .B(n6840), .C(n604), .Y(n3036) );
  NAND2X1 U1099 ( .A(\Mem[23][14] ), .B(n6842), .Y(n604) );
  OAI21X1 U1100 ( .A(n6576), .B(n6840), .C(n605), .Y(n3037) );
  NAND2X1 U1101 ( .A(\Mem[23][15] ), .B(n6841), .Y(n605) );
  OAI21X1 U1102 ( .A(n6571), .B(n6840), .C(n606), .Y(n3038) );
  NAND2X1 U1103 ( .A(\Mem[23][16] ), .B(n6842), .Y(n606) );
  OAI21X1 U1104 ( .A(n6566), .B(n6840), .C(n607), .Y(n3039) );
  NAND2X1 U1105 ( .A(\Mem[23][17] ), .B(n6841), .Y(n607) );
  OAI21X1 U1106 ( .A(n6561), .B(n6840), .C(n608), .Y(n3040) );
  NAND2X1 U1107 ( .A(\Mem[23][18] ), .B(n6841), .Y(n608) );
  OAI21X1 U1108 ( .A(n6555), .B(n6840), .C(n609), .Y(n3041) );
  NAND2X1 U1109 ( .A(\Mem[23][19] ), .B(n6841), .Y(n609) );
  OAI21X1 U1110 ( .A(n6545), .B(n6840), .C(n610), .Y(n3042) );
  NAND2X1 U1111 ( .A(\Mem[23][20] ), .B(n6841), .Y(n610) );
  OAI21X1 U1112 ( .A(n6540), .B(n6840), .C(n611), .Y(n3043) );
  NAND2X1 U1113 ( .A(\Mem[23][21] ), .B(n6841), .Y(n611) );
  OAI21X1 U1114 ( .A(n6535), .B(n6840), .C(n612), .Y(n3044) );
  NAND2X1 U1115 ( .A(\Mem[23][22] ), .B(n6842), .Y(n612) );
  OAI21X1 U1116 ( .A(n6530), .B(n6841), .C(n613), .Y(n3045) );
  NAND2X1 U1117 ( .A(\Mem[23][23] ), .B(n6841), .Y(n613) );
  OAI21X1 U1118 ( .A(n6525), .B(n6840), .C(n614), .Y(n3046) );
  NAND2X1 U1119 ( .A(\Mem[23][24] ), .B(n6842), .Y(n614) );
  OAI21X1 U1120 ( .A(n6520), .B(n6841), .C(n615), .Y(n3047) );
  NAND2X1 U1121 ( .A(\Mem[23][25] ), .B(n6842), .Y(n615) );
  OAI21X1 U1122 ( .A(n6515), .B(n6841), .C(n616), .Y(n3048) );
  NAND2X1 U1123 ( .A(\Mem[23][26] ), .B(n6842), .Y(n616) );
  OAI21X1 U1124 ( .A(n6510), .B(n6841), .C(n617), .Y(n3049) );
  NAND2X1 U1125 ( .A(\Mem[23][27] ), .B(n6842), .Y(n617) );
  OAI21X1 U1126 ( .A(n6505), .B(n6841), .C(n618), .Y(n3050) );
  NAND2X1 U1127 ( .A(\Mem[23][28] ), .B(n6842), .Y(n618) );
  OAI21X1 U1128 ( .A(n6500), .B(n6841), .C(n619), .Y(n3051) );
  NAND2X1 U1129 ( .A(\Mem[23][29] ), .B(n6842), .Y(n619) );
  OAI21X1 U1130 ( .A(n6490), .B(n6841), .C(n620), .Y(n3052) );
  NAND2X1 U1131 ( .A(\Mem[23][30] ), .B(n6843), .Y(n620) );
  OAI21X1 U1132 ( .A(n6485), .B(n6841), .C(n621), .Y(n3053) );
  NAND2X1 U1133 ( .A(\Mem[23][31] ), .B(n6843), .Y(n621) );
  NAND2X1 U1134 ( .A(n7006), .B(n7021), .Y(n589) );
  NAND3X1 U1136 ( .A(n81), .B(n7015), .C(ADDR_WR[4]), .Y(n622) );
  OAI21X1 U1137 ( .A(n6605), .B(n6835), .C(n625), .Y(n3054) );
  NAND2X1 U1138 ( .A(\Mem[24][0] ), .B(n6838), .Y(n625) );
  OAI21X1 U1139 ( .A(n6550), .B(n6834), .C(n626), .Y(n3055) );
  NAND2X1 U1140 ( .A(\Mem[24][1] ), .B(n6838), .Y(n626) );
  OAI21X1 U1141 ( .A(n6495), .B(n6834), .C(n627), .Y(n3056) );
  NAND2X1 U1142 ( .A(\Mem[24][2] ), .B(n6838), .Y(n627) );
  OAI21X1 U1143 ( .A(n6480), .B(n6834), .C(n628), .Y(n3057) );
  NAND2X1 U1144 ( .A(\Mem[24][3] ), .B(n6837), .Y(n628) );
  OAI21X1 U1145 ( .A(n6475), .B(n6834), .C(n629), .Y(n3058) );
  NAND2X1 U1146 ( .A(\Mem[24][4] ), .B(n6838), .Y(n629) );
  OAI21X1 U1147 ( .A(n6470), .B(n6834), .C(n630), .Y(n3059) );
  NAND2X1 U1148 ( .A(\Mem[24][5] ), .B(n6837), .Y(n630) );
  OAI21X1 U1149 ( .A(n6465), .B(n6834), .C(n631), .Y(n3060) );
  NAND2X1 U1150 ( .A(\Mem[24][6] ), .B(n6837), .Y(n631) );
  OAI21X1 U1151 ( .A(n6460), .B(n6834), .C(n632), .Y(n3061) );
  NAND2X1 U1152 ( .A(\Mem[24][7] ), .B(n6837), .Y(n632) );
  OAI21X1 U1153 ( .A(n6455), .B(n6834), .C(n633), .Y(n3062) );
  NAND2X1 U1154 ( .A(\Mem[24][8] ), .B(n6837), .Y(n633) );
  OAI21X1 U1155 ( .A(n6450), .B(n6834), .C(n634), .Y(n3063) );
  NAND2X1 U1156 ( .A(\Mem[24][9] ), .B(n6837), .Y(n634) );
  OAI21X1 U1157 ( .A(n6600), .B(n6834), .C(n635), .Y(n3064) );
  NAND2X1 U1158 ( .A(\Mem[24][10] ), .B(n6837), .Y(n635) );
  OAI21X1 U1159 ( .A(n6595), .B(n6834), .C(n636), .Y(n3065) );
  NAND2X1 U1160 ( .A(\Mem[24][11] ), .B(n6837), .Y(n636) );
  OAI21X1 U1161 ( .A(n6590), .B(n6834), .C(n637), .Y(n3066) );
  NAND2X1 U1162 ( .A(\Mem[24][12] ), .B(n6837), .Y(n637) );
  OAI21X1 U1163 ( .A(n6585), .B(n6835), .C(n638), .Y(n3067) );
  NAND2X1 U1164 ( .A(\Mem[24][13] ), .B(n6837), .Y(n638) );
  OAI21X1 U1165 ( .A(n6580), .B(n6835), .C(n639), .Y(n3068) );
  NAND2X1 U1166 ( .A(\Mem[24][14] ), .B(n6837), .Y(n639) );
  OAI21X1 U1167 ( .A(n6575), .B(n6835), .C(n640), .Y(n3069) );
  NAND2X1 U1168 ( .A(\Mem[24][15] ), .B(n6836), .Y(n640) );
  OAI21X1 U1169 ( .A(n6570), .B(n6835), .C(n641), .Y(n3070) );
  NAND2X1 U1170 ( .A(\Mem[24][16] ), .B(n6837), .Y(n641) );
  OAI21X1 U1171 ( .A(n6565), .B(n6835), .C(n642), .Y(n3071) );
  NAND2X1 U1172 ( .A(\Mem[24][17] ), .B(n6836), .Y(n642) );
  OAI21X1 U1173 ( .A(n6560), .B(n6835), .C(n643), .Y(n3072) );
  NAND2X1 U1174 ( .A(\Mem[24][18] ), .B(n6836), .Y(n643) );
  OAI21X1 U1175 ( .A(n6555), .B(n6835), .C(n644), .Y(n3073) );
  NAND2X1 U1176 ( .A(\Mem[24][19] ), .B(n6836), .Y(n644) );
  OAI21X1 U1177 ( .A(n6545), .B(n6835), .C(n645), .Y(n3074) );
  NAND2X1 U1178 ( .A(\Mem[24][20] ), .B(n6836), .Y(n645) );
  OAI21X1 U1179 ( .A(n6540), .B(n6835), .C(n646), .Y(n3075) );
  NAND2X1 U1180 ( .A(\Mem[24][21] ), .B(n6836), .Y(n646) );
  OAI21X1 U1181 ( .A(n6535), .B(n6835), .C(n647), .Y(n3076) );
  NAND2X1 U1182 ( .A(\Mem[24][22] ), .B(n6837), .Y(n647) );
  OAI21X1 U1183 ( .A(n6530), .B(n6836), .C(n648), .Y(n3077) );
  NAND2X1 U1184 ( .A(\Mem[24][23] ), .B(n6836), .Y(n648) );
  OAI21X1 U1185 ( .A(n6525), .B(n6835), .C(n649), .Y(n3078) );
  NAND2X1 U1186 ( .A(\Mem[24][24] ), .B(n6837), .Y(n649) );
  OAI21X1 U1187 ( .A(n6520), .B(n6836), .C(n650), .Y(n3079) );
  NAND2X1 U1188 ( .A(\Mem[24][25] ), .B(n6837), .Y(n650) );
  OAI21X1 U1189 ( .A(n6515), .B(n6836), .C(n651), .Y(n3080) );
  NAND2X1 U1190 ( .A(\Mem[24][26] ), .B(n6837), .Y(n651) );
  OAI21X1 U1191 ( .A(n6510), .B(n6836), .C(n652), .Y(n3081) );
  NAND2X1 U1192 ( .A(\Mem[24][27] ), .B(n6837), .Y(n652) );
  OAI21X1 U1193 ( .A(n6505), .B(n6836), .C(n653), .Y(n3082) );
  NAND2X1 U1194 ( .A(\Mem[24][28] ), .B(n6837), .Y(n653) );
  OAI21X1 U1195 ( .A(n6500), .B(n6836), .C(n654), .Y(n3083) );
  NAND2X1 U1196 ( .A(\Mem[24][29] ), .B(n6837), .Y(n654) );
  OAI21X1 U1197 ( .A(n6490), .B(n6836), .C(n655), .Y(n3084) );
  NAND2X1 U1198 ( .A(\Mem[24][30] ), .B(n6838), .Y(n655) );
  OAI21X1 U1199 ( .A(n6485), .B(n6836), .C(n656), .Y(n3085) );
  NAND2X1 U1200 ( .A(\Mem[24][31] ), .B(n6838), .Y(n656) );
  NAND2X1 U1201 ( .A(n7005), .B(n7016), .Y(n624) );
  OAI21X1 U1202 ( .A(n6605), .B(n6830), .C(n659), .Y(n3086) );
  NAND2X1 U1203 ( .A(\Mem[25][0] ), .B(n6833), .Y(n659) );
  OAI21X1 U1204 ( .A(n6550), .B(n6829), .C(n660), .Y(n3087) );
  NAND2X1 U1205 ( .A(\Mem[25][1] ), .B(n6833), .Y(n660) );
  OAI21X1 U1206 ( .A(n6495), .B(n6829), .C(n661), .Y(n3088) );
  NAND2X1 U1207 ( .A(\Mem[25][2] ), .B(n6833), .Y(n661) );
  OAI21X1 U1208 ( .A(n6480), .B(n6829), .C(n662), .Y(n3089) );
  NAND2X1 U1209 ( .A(\Mem[25][3] ), .B(n6832), .Y(n662) );
  OAI21X1 U1210 ( .A(n6475), .B(n6829), .C(n663), .Y(n3090) );
  NAND2X1 U1211 ( .A(\Mem[25][4] ), .B(n6833), .Y(n663) );
  OAI21X1 U1212 ( .A(n6470), .B(n6829), .C(n664), .Y(n3091) );
  NAND2X1 U1213 ( .A(\Mem[25][5] ), .B(n6832), .Y(n664) );
  OAI21X1 U1214 ( .A(n6465), .B(n6829), .C(n665), .Y(n3092) );
  NAND2X1 U1215 ( .A(\Mem[25][6] ), .B(n6832), .Y(n665) );
  OAI21X1 U1216 ( .A(n6460), .B(n6829), .C(n666), .Y(n3093) );
  NAND2X1 U1217 ( .A(\Mem[25][7] ), .B(n6832), .Y(n666) );
  OAI21X1 U1218 ( .A(n6455), .B(n6829), .C(n667), .Y(n3094) );
  NAND2X1 U1219 ( .A(\Mem[25][8] ), .B(n6832), .Y(n667) );
  OAI21X1 U1220 ( .A(n6450), .B(n6829), .C(n668), .Y(n3095) );
  NAND2X1 U1221 ( .A(\Mem[25][9] ), .B(n6832), .Y(n668) );
  OAI21X1 U1222 ( .A(n6600), .B(n6829), .C(n669), .Y(n3096) );
  NAND2X1 U1223 ( .A(\Mem[25][10] ), .B(n6832), .Y(n669) );
  OAI21X1 U1224 ( .A(n6595), .B(n6829), .C(n670), .Y(n3097) );
  NAND2X1 U1225 ( .A(\Mem[25][11] ), .B(n6832), .Y(n670) );
  OAI21X1 U1226 ( .A(n6590), .B(n6829), .C(n671), .Y(n3098) );
  NAND2X1 U1227 ( .A(\Mem[25][12] ), .B(n6832), .Y(n671) );
  OAI21X1 U1228 ( .A(n6585), .B(n6830), .C(n672), .Y(n3099) );
  NAND2X1 U1229 ( .A(\Mem[25][13] ), .B(n6832), .Y(n672) );
  OAI21X1 U1230 ( .A(n6580), .B(n6830), .C(n673), .Y(n3100) );
  NAND2X1 U1231 ( .A(\Mem[25][14] ), .B(n6832), .Y(n673) );
  OAI21X1 U1232 ( .A(n6575), .B(n6830), .C(n674), .Y(n3101) );
  NAND2X1 U1233 ( .A(\Mem[25][15] ), .B(n6831), .Y(n674) );
  OAI21X1 U1234 ( .A(n6570), .B(n6830), .C(n675), .Y(n3102) );
  NAND2X1 U1235 ( .A(\Mem[25][16] ), .B(n6832), .Y(n675) );
  OAI21X1 U1236 ( .A(n6565), .B(n6830), .C(n676), .Y(n3103) );
  NAND2X1 U1237 ( .A(\Mem[25][17] ), .B(n6831), .Y(n676) );
  OAI21X1 U1238 ( .A(n6560), .B(n6830), .C(n677), .Y(n3104) );
  NAND2X1 U1239 ( .A(\Mem[25][18] ), .B(n6831), .Y(n677) );
  OAI21X1 U1240 ( .A(n6555), .B(n6830), .C(n678), .Y(n3105) );
  NAND2X1 U1241 ( .A(\Mem[25][19] ), .B(n6831), .Y(n678) );
  OAI21X1 U1242 ( .A(n6545), .B(n6830), .C(n679), .Y(n3106) );
  NAND2X1 U1243 ( .A(\Mem[25][20] ), .B(n6831), .Y(n679) );
  OAI21X1 U1244 ( .A(n6540), .B(n6830), .C(n680), .Y(n3107) );
  NAND2X1 U1245 ( .A(\Mem[25][21] ), .B(n6831), .Y(n680) );
  OAI21X1 U1246 ( .A(n6535), .B(n6830), .C(n681), .Y(n3108) );
  NAND2X1 U1247 ( .A(\Mem[25][22] ), .B(n6832), .Y(n681) );
  OAI21X1 U1248 ( .A(n6530), .B(n6831), .C(n682), .Y(n3109) );
  NAND2X1 U1249 ( .A(\Mem[25][23] ), .B(n6831), .Y(n682) );
  OAI21X1 U1250 ( .A(n6525), .B(n6830), .C(n683), .Y(n3110) );
  NAND2X1 U1251 ( .A(\Mem[25][24] ), .B(n6832), .Y(n683) );
  OAI21X1 U1252 ( .A(n6520), .B(n6831), .C(n684), .Y(n3111) );
  NAND2X1 U1253 ( .A(\Mem[25][25] ), .B(n6832), .Y(n684) );
  OAI21X1 U1254 ( .A(n6515), .B(n6831), .C(n685), .Y(n3112) );
  NAND2X1 U1255 ( .A(\Mem[25][26] ), .B(n6832), .Y(n685) );
  OAI21X1 U1256 ( .A(n6510), .B(n6831), .C(n686), .Y(n3113) );
  NAND2X1 U1257 ( .A(\Mem[25][27] ), .B(n6832), .Y(n686) );
  OAI21X1 U1258 ( .A(n6505), .B(n6831), .C(n687), .Y(n3114) );
  NAND2X1 U1259 ( .A(\Mem[25][28] ), .B(n6832), .Y(n687) );
  OAI21X1 U1260 ( .A(n6500), .B(n6831), .C(n688), .Y(n3115) );
  NAND2X1 U1261 ( .A(\Mem[25][29] ), .B(n6832), .Y(n688) );
  OAI21X1 U1262 ( .A(n6490), .B(n6831), .C(n689), .Y(n3116) );
  NAND2X1 U1263 ( .A(\Mem[25][30] ), .B(n6833), .Y(n689) );
  OAI21X1 U1264 ( .A(n6485), .B(n6831), .C(n690), .Y(n3117) );
  NAND2X1 U1265 ( .A(\Mem[25][31] ), .B(n6833), .Y(n690) );
  NAND2X1 U1266 ( .A(n7005), .B(n7017), .Y(n658) );
  OAI21X1 U1267 ( .A(n6605), .B(n6825), .C(n692), .Y(n3118) );
  NAND2X1 U1268 ( .A(\Mem[26][0] ), .B(n6828), .Y(n692) );
  OAI21X1 U1269 ( .A(n6550), .B(n6824), .C(n693), .Y(n3119) );
  NAND2X1 U1270 ( .A(\Mem[26][1] ), .B(n6828), .Y(n693) );
  OAI21X1 U1271 ( .A(n6495), .B(n6824), .C(n694), .Y(n3120) );
  NAND2X1 U1272 ( .A(\Mem[26][2] ), .B(n6828), .Y(n694) );
  OAI21X1 U1273 ( .A(n6480), .B(n6824), .C(n695), .Y(n3121) );
  NAND2X1 U1274 ( .A(\Mem[26][3] ), .B(n6827), .Y(n695) );
  OAI21X1 U1275 ( .A(n6475), .B(n6824), .C(n696), .Y(n3122) );
  NAND2X1 U1276 ( .A(\Mem[26][4] ), .B(n6828), .Y(n696) );
  OAI21X1 U1277 ( .A(n6470), .B(n6824), .C(n697), .Y(n3123) );
  NAND2X1 U1278 ( .A(\Mem[26][5] ), .B(n6827), .Y(n697) );
  OAI21X1 U1279 ( .A(n6465), .B(n6824), .C(n698), .Y(n3124) );
  NAND2X1 U1280 ( .A(\Mem[26][6] ), .B(n6827), .Y(n698) );
  OAI21X1 U1281 ( .A(n6460), .B(n6824), .C(n699), .Y(n3125) );
  NAND2X1 U1282 ( .A(\Mem[26][7] ), .B(n6827), .Y(n699) );
  OAI21X1 U1283 ( .A(n6455), .B(n6824), .C(n700), .Y(n3126) );
  NAND2X1 U1284 ( .A(\Mem[26][8] ), .B(n6827), .Y(n700) );
  OAI21X1 U1285 ( .A(n6450), .B(n6824), .C(n701), .Y(n3127) );
  NAND2X1 U1286 ( .A(\Mem[26][9] ), .B(n6827), .Y(n701) );
  OAI21X1 U1287 ( .A(n6600), .B(n6824), .C(n702), .Y(n3128) );
  NAND2X1 U1288 ( .A(\Mem[26][10] ), .B(n6827), .Y(n702) );
  OAI21X1 U1289 ( .A(n6595), .B(n6824), .C(n703), .Y(n3129) );
  NAND2X1 U1290 ( .A(\Mem[26][11] ), .B(n6827), .Y(n703) );
  OAI21X1 U1291 ( .A(n6590), .B(n6824), .C(n704), .Y(n3130) );
  NAND2X1 U1292 ( .A(\Mem[26][12] ), .B(n6827), .Y(n704) );
  OAI21X1 U1293 ( .A(n6585), .B(n6825), .C(n705), .Y(n3131) );
  NAND2X1 U1294 ( .A(\Mem[26][13] ), .B(n6827), .Y(n705) );
  OAI21X1 U1295 ( .A(n6580), .B(n6825), .C(n706), .Y(n3132) );
  NAND2X1 U1296 ( .A(\Mem[26][14] ), .B(n6827), .Y(n706) );
  OAI21X1 U1297 ( .A(n6575), .B(n6825), .C(n707), .Y(n3133) );
  NAND2X1 U1298 ( .A(\Mem[26][15] ), .B(n6826), .Y(n707) );
  OAI21X1 U1299 ( .A(n6570), .B(n6825), .C(n708), .Y(n3134) );
  NAND2X1 U1300 ( .A(\Mem[26][16] ), .B(n6827), .Y(n708) );
  OAI21X1 U1301 ( .A(n6565), .B(n6825), .C(n709), .Y(n3135) );
  NAND2X1 U1302 ( .A(\Mem[26][17] ), .B(n6826), .Y(n709) );
  OAI21X1 U1303 ( .A(n6560), .B(n6825), .C(n710), .Y(n3136) );
  NAND2X1 U1304 ( .A(\Mem[26][18] ), .B(n6826), .Y(n710) );
  OAI21X1 U1305 ( .A(n6555), .B(n6825), .C(n711), .Y(n3137) );
  NAND2X1 U1306 ( .A(\Mem[26][19] ), .B(n6826), .Y(n711) );
  OAI21X1 U1307 ( .A(n6545), .B(n6825), .C(n712), .Y(n3138) );
  NAND2X1 U1308 ( .A(\Mem[26][20] ), .B(n6826), .Y(n712) );
  OAI21X1 U1309 ( .A(n6540), .B(n6825), .C(n713), .Y(n3139) );
  NAND2X1 U1310 ( .A(\Mem[26][21] ), .B(n6826), .Y(n713) );
  OAI21X1 U1311 ( .A(n6535), .B(n6825), .C(n714), .Y(n3140) );
  NAND2X1 U1312 ( .A(\Mem[26][22] ), .B(n6827), .Y(n714) );
  OAI21X1 U1313 ( .A(n6530), .B(n6826), .C(n715), .Y(n3141) );
  NAND2X1 U1314 ( .A(\Mem[26][23] ), .B(n6826), .Y(n715) );
  OAI21X1 U1315 ( .A(n6525), .B(n6825), .C(n716), .Y(n3142) );
  NAND2X1 U1316 ( .A(\Mem[26][24] ), .B(n6827), .Y(n716) );
  OAI21X1 U1317 ( .A(n6520), .B(n6826), .C(n717), .Y(n3143) );
  NAND2X1 U1318 ( .A(\Mem[26][25] ), .B(n6827), .Y(n717) );
  OAI21X1 U1319 ( .A(n6515), .B(n6826), .C(n718), .Y(n3144) );
  NAND2X1 U1320 ( .A(\Mem[26][26] ), .B(n6827), .Y(n718) );
  OAI21X1 U1321 ( .A(n6510), .B(n6826), .C(n719), .Y(n3145) );
  NAND2X1 U1322 ( .A(\Mem[26][27] ), .B(n6827), .Y(n719) );
  OAI21X1 U1323 ( .A(n6505), .B(n6826), .C(n720), .Y(n3146) );
  NAND2X1 U1324 ( .A(\Mem[26][28] ), .B(n6827), .Y(n720) );
  OAI21X1 U1325 ( .A(n6500), .B(n6826), .C(n721), .Y(n3147) );
  NAND2X1 U1326 ( .A(\Mem[26][29] ), .B(n6827), .Y(n721) );
  OAI21X1 U1327 ( .A(n6490), .B(n6826), .C(n722), .Y(n3148) );
  NAND2X1 U1328 ( .A(\Mem[26][30] ), .B(n6828), .Y(n722) );
  OAI21X1 U1329 ( .A(n6485), .B(n6826), .C(n723), .Y(n3149) );
  NAND2X1 U1330 ( .A(\Mem[26][31] ), .B(n6828), .Y(n723) );
  NAND2X1 U1331 ( .A(n7005), .B(n7018), .Y(n691) );
  OAI21X1 U1332 ( .A(n6605), .B(n6820), .C(n725), .Y(n3150) );
  NAND2X1 U1333 ( .A(\Mem[27][0] ), .B(n6823), .Y(n725) );
  OAI21X1 U1334 ( .A(n6550), .B(n6819), .C(n726), .Y(n3151) );
  NAND2X1 U1335 ( .A(\Mem[27][1] ), .B(n6823), .Y(n726) );
  OAI21X1 U1336 ( .A(n6495), .B(n6819), .C(n727), .Y(n3152) );
  NAND2X1 U1337 ( .A(\Mem[27][2] ), .B(n6823), .Y(n727) );
  OAI21X1 U1338 ( .A(n6480), .B(n6819), .C(n728), .Y(n3153) );
  NAND2X1 U1339 ( .A(\Mem[27][3] ), .B(n6822), .Y(n728) );
  OAI21X1 U1340 ( .A(n6475), .B(n6819), .C(n729), .Y(n3154) );
  NAND2X1 U1341 ( .A(\Mem[27][4] ), .B(n6823), .Y(n729) );
  OAI21X1 U1342 ( .A(n6470), .B(n6819), .C(n730), .Y(n3155) );
  NAND2X1 U1343 ( .A(\Mem[27][5] ), .B(n6822), .Y(n730) );
  OAI21X1 U1344 ( .A(n6465), .B(n6819), .C(n731), .Y(n3156) );
  NAND2X1 U1345 ( .A(\Mem[27][6] ), .B(n6822), .Y(n731) );
  OAI21X1 U1346 ( .A(n6460), .B(n6819), .C(n732), .Y(n3157) );
  NAND2X1 U1347 ( .A(\Mem[27][7] ), .B(n6822), .Y(n732) );
  OAI21X1 U1348 ( .A(n6455), .B(n6819), .C(n733), .Y(n3158) );
  NAND2X1 U1349 ( .A(\Mem[27][8] ), .B(n6822), .Y(n733) );
  OAI21X1 U1350 ( .A(n6450), .B(n6819), .C(n734), .Y(n3159) );
  NAND2X1 U1351 ( .A(\Mem[27][9] ), .B(n6822), .Y(n734) );
  OAI21X1 U1352 ( .A(n6600), .B(n6819), .C(n735), .Y(n3160) );
  NAND2X1 U1353 ( .A(\Mem[27][10] ), .B(n6822), .Y(n735) );
  OAI21X1 U1354 ( .A(n6595), .B(n6819), .C(n736), .Y(n3161) );
  NAND2X1 U1355 ( .A(\Mem[27][11] ), .B(n6822), .Y(n736) );
  OAI21X1 U1356 ( .A(n6590), .B(n6819), .C(n737), .Y(n3162) );
  NAND2X1 U1357 ( .A(\Mem[27][12] ), .B(n6822), .Y(n737) );
  OAI21X1 U1358 ( .A(n6585), .B(n6820), .C(n738), .Y(n3163) );
  NAND2X1 U1359 ( .A(\Mem[27][13] ), .B(n6822), .Y(n738) );
  OAI21X1 U1360 ( .A(n6580), .B(n6820), .C(n739), .Y(n3164) );
  NAND2X1 U1361 ( .A(\Mem[27][14] ), .B(n6822), .Y(n739) );
  OAI21X1 U1362 ( .A(n6575), .B(n6820), .C(n740), .Y(n3165) );
  NAND2X1 U1363 ( .A(\Mem[27][15] ), .B(n6821), .Y(n740) );
  OAI21X1 U1364 ( .A(n6570), .B(n6820), .C(n741), .Y(n3166) );
  NAND2X1 U1365 ( .A(\Mem[27][16] ), .B(n6822), .Y(n741) );
  OAI21X1 U1366 ( .A(n6565), .B(n6820), .C(n742), .Y(n3167) );
  NAND2X1 U1367 ( .A(\Mem[27][17] ), .B(n6821), .Y(n742) );
  OAI21X1 U1368 ( .A(n6560), .B(n6820), .C(n743), .Y(n3168) );
  NAND2X1 U1369 ( .A(\Mem[27][18] ), .B(n6821), .Y(n743) );
  OAI21X1 U1370 ( .A(n6555), .B(n6820), .C(n744), .Y(n3169) );
  NAND2X1 U1371 ( .A(\Mem[27][19] ), .B(n6821), .Y(n744) );
  OAI21X1 U1372 ( .A(n6545), .B(n6820), .C(n745), .Y(n3170) );
  NAND2X1 U1373 ( .A(\Mem[27][20] ), .B(n6821), .Y(n745) );
  OAI21X1 U1374 ( .A(n6540), .B(n6820), .C(n746), .Y(n3171) );
  NAND2X1 U1375 ( .A(\Mem[27][21] ), .B(n6821), .Y(n746) );
  OAI21X1 U1376 ( .A(n6535), .B(n6820), .C(n747), .Y(n3172) );
  NAND2X1 U1377 ( .A(\Mem[27][22] ), .B(n6822), .Y(n747) );
  OAI21X1 U1378 ( .A(n6530), .B(n6821), .C(n748), .Y(n3173) );
  NAND2X1 U1379 ( .A(\Mem[27][23] ), .B(n6821), .Y(n748) );
  OAI21X1 U1380 ( .A(n6525), .B(n6820), .C(n749), .Y(n3174) );
  NAND2X1 U1381 ( .A(\Mem[27][24] ), .B(n6822), .Y(n749) );
  OAI21X1 U1382 ( .A(n6520), .B(n6821), .C(n750), .Y(n3175) );
  NAND2X1 U1383 ( .A(\Mem[27][25] ), .B(n6822), .Y(n750) );
  OAI21X1 U1384 ( .A(n6515), .B(n6821), .C(n751), .Y(n3176) );
  NAND2X1 U1385 ( .A(\Mem[27][26] ), .B(n6822), .Y(n751) );
  OAI21X1 U1386 ( .A(n6510), .B(n6821), .C(n752), .Y(n3177) );
  NAND2X1 U1387 ( .A(\Mem[27][27] ), .B(n6822), .Y(n752) );
  OAI21X1 U1388 ( .A(n6505), .B(n6821), .C(n753), .Y(n3178) );
  NAND2X1 U1389 ( .A(\Mem[27][28] ), .B(n6822), .Y(n753) );
  OAI21X1 U1390 ( .A(n6500), .B(n6821), .C(n754), .Y(n3179) );
  NAND2X1 U1391 ( .A(\Mem[27][29] ), .B(n6822), .Y(n754) );
  OAI21X1 U1392 ( .A(n6490), .B(n6821), .C(n755), .Y(n3180) );
  NAND2X1 U1393 ( .A(\Mem[27][30] ), .B(n6823), .Y(n755) );
  OAI21X1 U1394 ( .A(n6485), .B(n6821), .C(n756), .Y(n3181) );
  NAND2X1 U1395 ( .A(\Mem[27][31] ), .B(n6823), .Y(n756) );
  NAND2X1 U1396 ( .A(n7005), .B(n7019), .Y(n724) );
  OAI21X1 U1397 ( .A(n6605), .B(n6815), .C(n758), .Y(n3182) );
  NAND2X1 U1398 ( .A(\Mem[28][0] ), .B(n6818), .Y(n758) );
  OAI21X1 U1399 ( .A(n6550), .B(n6814), .C(n759), .Y(n3183) );
  NAND2X1 U1400 ( .A(\Mem[28][1] ), .B(n6818), .Y(n759) );
  OAI21X1 U1401 ( .A(n6495), .B(n6814), .C(n760), .Y(n3184) );
  NAND2X1 U1402 ( .A(\Mem[28][2] ), .B(n6818), .Y(n760) );
  OAI21X1 U1403 ( .A(n6480), .B(n6814), .C(n761), .Y(n3185) );
  NAND2X1 U1404 ( .A(\Mem[28][3] ), .B(n6817), .Y(n761) );
  OAI21X1 U1405 ( .A(n6475), .B(n6814), .C(n762), .Y(n3186) );
  NAND2X1 U1406 ( .A(\Mem[28][4] ), .B(n6818), .Y(n762) );
  OAI21X1 U1407 ( .A(n6470), .B(n6814), .C(n763), .Y(n3187) );
  NAND2X1 U1408 ( .A(\Mem[28][5] ), .B(n6817), .Y(n763) );
  OAI21X1 U1409 ( .A(n6465), .B(n6814), .C(n764), .Y(n3188) );
  NAND2X1 U1410 ( .A(\Mem[28][6] ), .B(n6817), .Y(n764) );
  OAI21X1 U1411 ( .A(n6460), .B(n6814), .C(n765), .Y(n3189) );
  NAND2X1 U1412 ( .A(\Mem[28][7] ), .B(n6817), .Y(n765) );
  OAI21X1 U1413 ( .A(n6455), .B(n6814), .C(n766), .Y(n3190) );
  NAND2X1 U1414 ( .A(\Mem[28][8] ), .B(n6817), .Y(n766) );
  OAI21X1 U1415 ( .A(n6450), .B(n6814), .C(n767), .Y(n3191) );
  NAND2X1 U1416 ( .A(\Mem[28][9] ), .B(n6817), .Y(n767) );
  OAI21X1 U1417 ( .A(n6600), .B(n6814), .C(n768), .Y(n3192) );
  NAND2X1 U1418 ( .A(\Mem[28][10] ), .B(n6817), .Y(n768) );
  OAI21X1 U1419 ( .A(n6595), .B(n6814), .C(n769), .Y(n3193) );
  NAND2X1 U1420 ( .A(\Mem[28][11] ), .B(n6817), .Y(n769) );
  OAI21X1 U1421 ( .A(n6590), .B(n6814), .C(n770), .Y(n3194) );
  NAND2X1 U1422 ( .A(\Mem[28][12] ), .B(n6817), .Y(n770) );
  OAI21X1 U1423 ( .A(n6585), .B(n6815), .C(n771), .Y(n3195) );
  NAND2X1 U1424 ( .A(\Mem[28][13] ), .B(n6817), .Y(n771) );
  OAI21X1 U1425 ( .A(n6580), .B(n6815), .C(n772), .Y(n3196) );
  NAND2X1 U1426 ( .A(\Mem[28][14] ), .B(n6817), .Y(n772) );
  OAI21X1 U1427 ( .A(n6575), .B(n6815), .C(n773), .Y(n3197) );
  NAND2X1 U1428 ( .A(\Mem[28][15] ), .B(n6816), .Y(n773) );
  OAI21X1 U1429 ( .A(n6570), .B(n6815), .C(n774), .Y(n3198) );
  NAND2X1 U1430 ( .A(\Mem[28][16] ), .B(n6817), .Y(n774) );
  OAI21X1 U1431 ( .A(n6565), .B(n6815), .C(n775), .Y(n3199) );
  NAND2X1 U1432 ( .A(\Mem[28][17] ), .B(n6816), .Y(n775) );
  OAI21X1 U1433 ( .A(n6560), .B(n6815), .C(n776), .Y(n3200) );
  NAND2X1 U1434 ( .A(\Mem[28][18] ), .B(n6816), .Y(n776) );
  OAI21X1 U1435 ( .A(n6555), .B(n6815), .C(n777), .Y(n3201) );
  NAND2X1 U1436 ( .A(\Mem[28][19] ), .B(n6816), .Y(n777) );
  OAI21X1 U1437 ( .A(n6545), .B(n6815), .C(n778), .Y(n3202) );
  NAND2X1 U1438 ( .A(\Mem[28][20] ), .B(n6816), .Y(n778) );
  OAI21X1 U1439 ( .A(n6540), .B(n6815), .C(n779), .Y(n3203) );
  NAND2X1 U1440 ( .A(\Mem[28][21] ), .B(n6816), .Y(n779) );
  OAI21X1 U1441 ( .A(n6535), .B(n6815), .C(n780), .Y(n3204) );
  NAND2X1 U1442 ( .A(\Mem[28][22] ), .B(n6817), .Y(n780) );
  OAI21X1 U1443 ( .A(n6530), .B(n6816), .C(n781), .Y(n3205) );
  NAND2X1 U1444 ( .A(\Mem[28][23] ), .B(n6816), .Y(n781) );
  OAI21X1 U1445 ( .A(n6525), .B(n6815), .C(n782), .Y(n3206) );
  NAND2X1 U1446 ( .A(\Mem[28][24] ), .B(n6817), .Y(n782) );
  OAI21X1 U1447 ( .A(n6520), .B(n6816), .C(n783), .Y(n3207) );
  NAND2X1 U1448 ( .A(\Mem[28][25] ), .B(n6817), .Y(n783) );
  OAI21X1 U1449 ( .A(n6515), .B(n6816), .C(n784), .Y(n3208) );
  NAND2X1 U1450 ( .A(\Mem[28][26] ), .B(n6817), .Y(n784) );
  OAI21X1 U1451 ( .A(n6510), .B(n6816), .C(n785), .Y(n3209) );
  NAND2X1 U1452 ( .A(\Mem[28][27] ), .B(n6817), .Y(n785) );
  OAI21X1 U1453 ( .A(n6505), .B(n6816), .C(n786), .Y(n3210) );
  NAND2X1 U1454 ( .A(\Mem[28][28] ), .B(n6817), .Y(n786) );
  OAI21X1 U1455 ( .A(n6500), .B(n6816), .C(n787), .Y(n3211) );
  NAND2X1 U1456 ( .A(\Mem[28][29] ), .B(n6817), .Y(n787) );
  OAI21X1 U1457 ( .A(n6490), .B(n6816), .C(n788), .Y(n3212) );
  NAND2X1 U1458 ( .A(\Mem[28][30] ), .B(n6818), .Y(n788) );
  OAI21X1 U1459 ( .A(n6485), .B(n6816), .C(n789), .Y(n3213) );
  NAND2X1 U1460 ( .A(\Mem[28][31] ), .B(n6818), .Y(n789) );
  NAND2X1 U1461 ( .A(n7005), .B(n7022), .Y(n757) );
  OAI21X1 U1462 ( .A(n6605), .B(n6810), .C(n791), .Y(n3214) );
  NAND2X1 U1463 ( .A(\Mem[29][0] ), .B(n6813), .Y(n791) );
  OAI21X1 U1464 ( .A(n6550), .B(n6809), .C(n792), .Y(n3215) );
  NAND2X1 U1465 ( .A(\Mem[29][1] ), .B(n6813), .Y(n792) );
  OAI21X1 U1466 ( .A(n6495), .B(n6809), .C(n793), .Y(n3216) );
  NAND2X1 U1467 ( .A(\Mem[29][2] ), .B(n6813), .Y(n793) );
  OAI21X1 U1468 ( .A(n6480), .B(n6809), .C(n794), .Y(n3217) );
  NAND2X1 U1469 ( .A(\Mem[29][3] ), .B(n6812), .Y(n794) );
  OAI21X1 U1470 ( .A(n6475), .B(n6809), .C(n795), .Y(n3218) );
  NAND2X1 U1471 ( .A(\Mem[29][4] ), .B(n6813), .Y(n795) );
  OAI21X1 U1472 ( .A(n6470), .B(n6809), .C(n796), .Y(n3219) );
  NAND2X1 U1473 ( .A(\Mem[29][5] ), .B(n6812), .Y(n796) );
  OAI21X1 U1474 ( .A(n6465), .B(n6809), .C(n797), .Y(n3220) );
  NAND2X1 U1475 ( .A(\Mem[29][6] ), .B(n6812), .Y(n797) );
  OAI21X1 U1476 ( .A(n6460), .B(n6809), .C(n798), .Y(n3221) );
  NAND2X1 U1477 ( .A(\Mem[29][7] ), .B(n6812), .Y(n798) );
  OAI21X1 U1478 ( .A(n6455), .B(n6809), .C(n799), .Y(n3222) );
  NAND2X1 U1479 ( .A(\Mem[29][8] ), .B(n6812), .Y(n799) );
  OAI21X1 U1480 ( .A(n6450), .B(n6809), .C(n800), .Y(n3223) );
  NAND2X1 U1481 ( .A(\Mem[29][9] ), .B(n6812), .Y(n800) );
  OAI21X1 U1482 ( .A(n6600), .B(n6809), .C(n801), .Y(n3224) );
  NAND2X1 U1483 ( .A(\Mem[29][10] ), .B(n6812), .Y(n801) );
  OAI21X1 U1484 ( .A(n6595), .B(n6809), .C(n802), .Y(n3225) );
  NAND2X1 U1485 ( .A(\Mem[29][11] ), .B(n6812), .Y(n802) );
  OAI21X1 U1486 ( .A(n6590), .B(n6809), .C(n803), .Y(n3226) );
  NAND2X1 U1487 ( .A(\Mem[29][12] ), .B(n6812), .Y(n803) );
  OAI21X1 U1488 ( .A(n6585), .B(n6810), .C(n804), .Y(n3227) );
  NAND2X1 U1489 ( .A(\Mem[29][13] ), .B(n6812), .Y(n804) );
  OAI21X1 U1490 ( .A(n6580), .B(n6810), .C(n805), .Y(n3228) );
  NAND2X1 U1491 ( .A(\Mem[29][14] ), .B(n6812), .Y(n805) );
  OAI21X1 U1492 ( .A(n6575), .B(n6810), .C(n806), .Y(n3229) );
  NAND2X1 U1493 ( .A(\Mem[29][15] ), .B(n6811), .Y(n806) );
  OAI21X1 U1494 ( .A(n6570), .B(n6810), .C(n807), .Y(n3230) );
  NAND2X1 U1495 ( .A(\Mem[29][16] ), .B(n6812), .Y(n807) );
  OAI21X1 U1496 ( .A(n6565), .B(n6810), .C(n808), .Y(n3231) );
  NAND2X1 U1497 ( .A(\Mem[29][17] ), .B(n6811), .Y(n808) );
  OAI21X1 U1498 ( .A(n6560), .B(n6810), .C(n809), .Y(n3232) );
  NAND2X1 U1499 ( .A(\Mem[29][18] ), .B(n6811), .Y(n809) );
  OAI21X1 U1500 ( .A(n6555), .B(n6810), .C(n810), .Y(n3233) );
  NAND2X1 U1501 ( .A(\Mem[29][19] ), .B(n6811), .Y(n810) );
  OAI21X1 U1502 ( .A(n6545), .B(n6810), .C(n811), .Y(n3234) );
  NAND2X1 U1503 ( .A(\Mem[29][20] ), .B(n6811), .Y(n811) );
  OAI21X1 U1504 ( .A(n6540), .B(n6810), .C(n812), .Y(n3235) );
  NAND2X1 U1505 ( .A(\Mem[29][21] ), .B(n6811), .Y(n812) );
  OAI21X1 U1506 ( .A(n6535), .B(n6810), .C(n813), .Y(n3236) );
  NAND2X1 U1507 ( .A(\Mem[29][22] ), .B(n6812), .Y(n813) );
  OAI21X1 U1508 ( .A(n6530), .B(n6811), .C(n814), .Y(n3237) );
  NAND2X1 U1509 ( .A(\Mem[29][23] ), .B(n6811), .Y(n814) );
  OAI21X1 U1510 ( .A(n6525), .B(n6810), .C(n815), .Y(n3238) );
  NAND2X1 U1511 ( .A(\Mem[29][24] ), .B(n6812), .Y(n815) );
  OAI21X1 U1512 ( .A(n6520), .B(n6811), .C(n816), .Y(n3239) );
  NAND2X1 U1513 ( .A(\Mem[29][25] ), .B(n6812), .Y(n816) );
  OAI21X1 U1514 ( .A(n6515), .B(n6811), .C(n817), .Y(n3240) );
  NAND2X1 U1515 ( .A(\Mem[29][26] ), .B(n6812), .Y(n817) );
  OAI21X1 U1516 ( .A(n6510), .B(n6811), .C(n818), .Y(n3241) );
  NAND2X1 U1517 ( .A(\Mem[29][27] ), .B(n6812), .Y(n818) );
  OAI21X1 U1518 ( .A(n6505), .B(n6811), .C(n819), .Y(n3242) );
  NAND2X1 U1519 ( .A(\Mem[29][28] ), .B(n6812), .Y(n819) );
  OAI21X1 U1520 ( .A(n6500), .B(n6811), .C(n820), .Y(n3243) );
  NAND2X1 U1521 ( .A(\Mem[29][29] ), .B(n6812), .Y(n820) );
  OAI21X1 U1522 ( .A(n6490), .B(n6811), .C(n821), .Y(n3244) );
  NAND2X1 U1523 ( .A(\Mem[29][30] ), .B(n6813), .Y(n821) );
  OAI21X1 U1524 ( .A(n6485), .B(n6811), .C(n822), .Y(n3245) );
  NAND2X1 U1525 ( .A(\Mem[29][31] ), .B(n6813), .Y(n822) );
  NAND2X1 U1526 ( .A(n7005), .B(n7023), .Y(n790) );
  OAI21X1 U1527 ( .A(n6605), .B(n6805), .C(n824), .Y(n3246) );
  NAND2X1 U1528 ( .A(\Mem[30][0] ), .B(n6808), .Y(n824) );
  OAI21X1 U1529 ( .A(n6550), .B(n6804), .C(n825), .Y(n3247) );
  NAND2X1 U1530 ( .A(\Mem[30][1] ), .B(n6808), .Y(n825) );
  OAI21X1 U1531 ( .A(n6495), .B(n6804), .C(n826), .Y(n3248) );
  NAND2X1 U1532 ( .A(\Mem[30][2] ), .B(n6808), .Y(n826) );
  OAI21X1 U1533 ( .A(n6480), .B(n6804), .C(n827), .Y(n3249) );
  NAND2X1 U1534 ( .A(\Mem[30][3] ), .B(n6807), .Y(n827) );
  OAI21X1 U1535 ( .A(n6475), .B(n6804), .C(n828), .Y(n3250) );
  NAND2X1 U1536 ( .A(\Mem[30][4] ), .B(n6808), .Y(n828) );
  OAI21X1 U1537 ( .A(n6470), .B(n6804), .C(n829), .Y(n3251) );
  NAND2X1 U1538 ( .A(\Mem[30][5] ), .B(n6807), .Y(n829) );
  OAI21X1 U1539 ( .A(n6465), .B(n6804), .C(n830), .Y(n3252) );
  NAND2X1 U1540 ( .A(\Mem[30][6] ), .B(n6807), .Y(n830) );
  OAI21X1 U1541 ( .A(n6460), .B(n6804), .C(n831), .Y(n3253) );
  NAND2X1 U1542 ( .A(\Mem[30][7] ), .B(n6807), .Y(n831) );
  OAI21X1 U1543 ( .A(n6455), .B(n6804), .C(n832), .Y(n3254) );
  NAND2X1 U1544 ( .A(\Mem[30][8] ), .B(n6807), .Y(n832) );
  OAI21X1 U1545 ( .A(n6450), .B(n6804), .C(n833), .Y(n3255) );
  NAND2X1 U1546 ( .A(\Mem[30][9] ), .B(n6807), .Y(n833) );
  OAI21X1 U1547 ( .A(n6600), .B(n6804), .C(n834), .Y(n3256) );
  NAND2X1 U1548 ( .A(\Mem[30][10] ), .B(n6807), .Y(n834) );
  OAI21X1 U1549 ( .A(n6595), .B(n6804), .C(n835), .Y(n3257) );
  NAND2X1 U1550 ( .A(\Mem[30][11] ), .B(n6807), .Y(n835) );
  OAI21X1 U1551 ( .A(n6590), .B(n6804), .C(n836), .Y(n3258) );
  NAND2X1 U1552 ( .A(\Mem[30][12] ), .B(n6807), .Y(n836) );
  OAI21X1 U1553 ( .A(n6585), .B(n6805), .C(n837), .Y(n3259) );
  NAND2X1 U1554 ( .A(\Mem[30][13] ), .B(n6807), .Y(n837) );
  OAI21X1 U1555 ( .A(n6580), .B(n6805), .C(n838), .Y(n3260) );
  NAND2X1 U1556 ( .A(\Mem[30][14] ), .B(n6807), .Y(n838) );
  OAI21X1 U1557 ( .A(n6575), .B(n6805), .C(n839), .Y(n3261) );
  NAND2X1 U1558 ( .A(\Mem[30][15] ), .B(n6806), .Y(n839) );
  OAI21X1 U1559 ( .A(n6570), .B(n6805), .C(n840), .Y(n3262) );
  NAND2X1 U1560 ( .A(\Mem[30][16] ), .B(n6807), .Y(n840) );
  OAI21X1 U1561 ( .A(n6565), .B(n6805), .C(n841), .Y(n3263) );
  NAND2X1 U1562 ( .A(\Mem[30][17] ), .B(n6806), .Y(n841) );
  OAI21X1 U1563 ( .A(n6560), .B(n6805), .C(n842), .Y(n3264) );
  NAND2X1 U1564 ( .A(\Mem[30][18] ), .B(n6806), .Y(n842) );
  OAI21X1 U1565 ( .A(n6555), .B(n6805), .C(n843), .Y(n3265) );
  NAND2X1 U1566 ( .A(\Mem[30][19] ), .B(n6806), .Y(n843) );
  OAI21X1 U1567 ( .A(n6545), .B(n6805), .C(n844), .Y(n3266) );
  NAND2X1 U1568 ( .A(\Mem[30][20] ), .B(n6806), .Y(n844) );
  OAI21X1 U1569 ( .A(n6540), .B(n6805), .C(n845), .Y(n3267) );
  NAND2X1 U1570 ( .A(\Mem[30][21] ), .B(n6806), .Y(n845) );
  OAI21X1 U1571 ( .A(n6535), .B(n6805), .C(n846), .Y(n3268) );
  NAND2X1 U1572 ( .A(\Mem[30][22] ), .B(n6807), .Y(n846) );
  OAI21X1 U1573 ( .A(n6530), .B(n6806), .C(n847), .Y(n3269) );
  NAND2X1 U1574 ( .A(\Mem[30][23] ), .B(n6806), .Y(n847) );
  OAI21X1 U1575 ( .A(n6525), .B(n6805), .C(n848), .Y(n3270) );
  NAND2X1 U1576 ( .A(\Mem[30][24] ), .B(n6807), .Y(n848) );
  OAI21X1 U1577 ( .A(n6520), .B(n6806), .C(n849), .Y(n3271) );
  NAND2X1 U1578 ( .A(\Mem[30][25] ), .B(n6807), .Y(n849) );
  OAI21X1 U1579 ( .A(n6515), .B(n6806), .C(n850), .Y(n3272) );
  NAND2X1 U1580 ( .A(\Mem[30][26] ), .B(n6807), .Y(n850) );
  OAI21X1 U1581 ( .A(n6510), .B(n6806), .C(n851), .Y(n3273) );
  NAND2X1 U1582 ( .A(\Mem[30][27] ), .B(n6807), .Y(n851) );
  OAI21X1 U1583 ( .A(n6505), .B(n6806), .C(n852), .Y(n3274) );
  NAND2X1 U1584 ( .A(\Mem[30][28] ), .B(n6807), .Y(n852) );
  OAI21X1 U1585 ( .A(n6500), .B(n6806), .C(n853), .Y(n3275) );
  NAND2X1 U1586 ( .A(\Mem[30][29] ), .B(n6807), .Y(n853) );
  OAI21X1 U1587 ( .A(n6490), .B(n6806), .C(n854), .Y(n3276) );
  NAND2X1 U1588 ( .A(\Mem[30][30] ), .B(n6808), .Y(n854) );
  OAI21X1 U1589 ( .A(n6485), .B(n6806), .C(n855), .Y(n3277) );
  NAND2X1 U1590 ( .A(\Mem[30][31] ), .B(n6808), .Y(n855) );
  NAND2X1 U1591 ( .A(n7005), .B(n7024), .Y(n823) );
  OAI21X1 U1592 ( .A(n6605), .B(n6800), .C(n857), .Y(n3278) );
  NAND2X1 U1593 ( .A(\Mem[31][0] ), .B(n6803), .Y(n857) );
  OAI21X1 U1594 ( .A(n6550), .B(n6799), .C(n858), .Y(n3279) );
  NAND2X1 U1595 ( .A(\Mem[31][1] ), .B(n6803), .Y(n858) );
  OAI21X1 U1596 ( .A(n6495), .B(n6799), .C(n859), .Y(n3280) );
  NAND2X1 U1597 ( .A(\Mem[31][2] ), .B(n6803), .Y(n859) );
  OAI21X1 U1598 ( .A(n6480), .B(n6799), .C(n860), .Y(n3281) );
  NAND2X1 U1599 ( .A(\Mem[31][3] ), .B(n6802), .Y(n860) );
  OAI21X1 U1600 ( .A(n6475), .B(n6799), .C(n861), .Y(n3282) );
  NAND2X1 U1601 ( .A(\Mem[31][4] ), .B(n6803), .Y(n861) );
  OAI21X1 U1602 ( .A(n6470), .B(n6799), .C(n862), .Y(n3283) );
  NAND2X1 U1603 ( .A(\Mem[31][5] ), .B(n6802), .Y(n862) );
  OAI21X1 U1604 ( .A(n6465), .B(n6799), .C(n863), .Y(n3284) );
  NAND2X1 U1605 ( .A(\Mem[31][6] ), .B(n6802), .Y(n863) );
  OAI21X1 U1606 ( .A(n6460), .B(n6799), .C(n864), .Y(n3285) );
  NAND2X1 U1607 ( .A(\Mem[31][7] ), .B(n6802), .Y(n864) );
  OAI21X1 U1608 ( .A(n6455), .B(n6799), .C(n865), .Y(n3286) );
  NAND2X1 U1609 ( .A(\Mem[31][8] ), .B(n6802), .Y(n865) );
  OAI21X1 U1610 ( .A(n6450), .B(n6799), .C(n866), .Y(n3287) );
  NAND2X1 U1611 ( .A(\Mem[31][9] ), .B(n6802), .Y(n866) );
  OAI21X1 U1612 ( .A(n6600), .B(n6799), .C(n867), .Y(n3288) );
  NAND2X1 U1613 ( .A(\Mem[31][10] ), .B(n6802), .Y(n867) );
  OAI21X1 U1614 ( .A(n6595), .B(n6799), .C(n868), .Y(n3289) );
  NAND2X1 U1615 ( .A(\Mem[31][11] ), .B(n6802), .Y(n868) );
  OAI21X1 U1616 ( .A(n6590), .B(n6799), .C(n869), .Y(n3290) );
  NAND2X1 U1617 ( .A(\Mem[31][12] ), .B(n6802), .Y(n869) );
  OAI21X1 U1618 ( .A(n6585), .B(n6800), .C(n870), .Y(n3291) );
  NAND2X1 U1619 ( .A(\Mem[31][13] ), .B(n6802), .Y(n870) );
  OAI21X1 U1620 ( .A(n6580), .B(n6800), .C(n871), .Y(n3292) );
  NAND2X1 U1621 ( .A(\Mem[31][14] ), .B(n6802), .Y(n871) );
  OAI21X1 U1622 ( .A(n6575), .B(n6800), .C(n872), .Y(n3293) );
  NAND2X1 U1623 ( .A(\Mem[31][15] ), .B(n6801), .Y(n872) );
  OAI21X1 U1624 ( .A(n6570), .B(n6800), .C(n873), .Y(n3294) );
  NAND2X1 U1625 ( .A(\Mem[31][16] ), .B(n6802), .Y(n873) );
  OAI21X1 U1626 ( .A(n6565), .B(n6800), .C(n874), .Y(n3295) );
  NAND2X1 U1627 ( .A(\Mem[31][17] ), .B(n6801), .Y(n874) );
  OAI21X1 U1628 ( .A(n6560), .B(n6800), .C(n875), .Y(n3296) );
  NAND2X1 U1629 ( .A(\Mem[31][18] ), .B(n6801), .Y(n875) );
  OAI21X1 U1630 ( .A(n6555), .B(n6800), .C(n876), .Y(n3297) );
  NAND2X1 U1631 ( .A(\Mem[31][19] ), .B(n6801), .Y(n876) );
  OAI21X1 U1632 ( .A(n6545), .B(n6800), .C(n877), .Y(n3298) );
  NAND2X1 U1633 ( .A(\Mem[31][20] ), .B(n6801), .Y(n877) );
  OAI21X1 U1634 ( .A(n6540), .B(n6800), .C(n878), .Y(n3299) );
  NAND2X1 U1635 ( .A(\Mem[31][21] ), .B(n6801), .Y(n878) );
  OAI21X1 U1636 ( .A(n6535), .B(n6800), .C(n879), .Y(n3300) );
  NAND2X1 U1637 ( .A(\Mem[31][22] ), .B(n6802), .Y(n879) );
  OAI21X1 U1638 ( .A(n6530), .B(n6801), .C(n880), .Y(n3301) );
  NAND2X1 U1639 ( .A(\Mem[31][23] ), .B(n6801), .Y(n880) );
  OAI21X1 U1640 ( .A(n6525), .B(n6800), .C(n881), .Y(n3302) );
  NAND2X1 U1641 ( .A(\Mem[31][24] ), .B(n6802), .Y(n881) );
  OAI21X1 U1642 ( .A(n6520), .B(n6801), .C(n882), .Y(n3303) );
  NAND2X1 U1643 ( .A(\Mem[31][25] ), .B(n6802), .Y(n882) );
  OAI21X1 U1644 ( .A(n6515), .B(n6801), .C(n883), .Y(n3304) );
  NAND2X1 U1645 ( .A(\Mem[31][26] ), .B(n6802), .Y(n883) );
  OAI21X1 U1646 ( .A(n6510), .B(n6801), .C(n884), .Y(n3305) );
  NAND2X1 U1647 ( .A(\Mem[31][27] ), .B(n6802), .Y(n884) );
  OAI21X1 U1648 ( .A(n6505), .B(n6801), .C(n885), .Y(n3306) );
  NAND2X1 U1649 ( .A(\Mem[31][28] ), .B(n6802), .Y(n885) );
  OAI21X1 U1650 ( .A(n6500), .B(n6801), .C(n886), .Y(n3307) );
  NAND2X1 U1651 ( .A(\Mem[31][29] ), .B(n6802), .Y(n886) );
  OAI21X1 U1652 ( .A(n6490), .B(n6801), .C(n887), .Y(n3308) );
  NAND2X1 U1653 ( .A(\Mem[31][30] ), .B(n6803), .Y(n887) );
  OAI21X1 U1654 ( .A(n6485), .B(n6801), .C(n888), .Y(n3309) );
  NAND2X1 U1655 ( .A(\Mem[31][31] ), .B(n6803), .Y(n888) );
  NAND2X1 U1656 ( .A(n7005), .B(n7021), .Y(n856) );
  NAND3X1 U1658 ( .A(ADDR_WR[3]), .B(n355), .C(ADDR_WR[4]), .Y(n889) );
  OAI21X1 U1659 ( .A(n6606), .B(n6795), .C(n891), .Y(n3310) );
  NAND2X1 U1660 ( .A(\Mem[32][0] ), .B(n6798), .Y(n891) );
  OAI21X1 U1661 ( .A(n6551), .B(n6794), .C(n892), .Y(n3311) );
  NAND2X1 U1662 ( .A(\Mem[32][1] ), .B(n6798), .Y(n892) );
  OAI21X1 U1663 ( .A(n6496), .B(n6794), .C(n893), .Y(n3312) );
  NAND2X1 U1664 ( .A(\Mem[32][2] ), .B(n6798), .Y(n893) );
  OAI21X1 U1665 ( .A(n6481), .B(n6794), .C(n894), .Y(n3313) );
  NAND2X1 U1666 ( .A(\Mem[32][3] ), .B(n6797), .Y(n894) );
  OAI21X1 U1667 ( .A(n6476), .B(n6794), .C(n895), .Y(n3314) );
  NAND2X1 U1668 ( .A(\Mem[32][4] ), .B(n6798), .Y(n895) );
  OAI21X1 U1669 ( .A(n6471), .B(n6794), .C(n896), .Y(n3315) );
  NAND2X1 U1670 ( .A(\Mem[32][5] ), .B(n6797), .Y(n896) );
  OAI21X1 U1671 ( .A(n6466), .B(n6794), .C(n897), .Y(n3316) );
  NAND2X1 U1672 ( .A(\Mem[32][6] ), .B(n6797), .Y(n897) );
  OAI21X1 U1673 ( .A(n6461), .B(n6794), .C(n898), .Y(n3317) );
  NAND2X1 U1674 ( .A(\Mem[32][7] ), .B(n6797), .Y(n898) );
  OAI21X1 U1675 ( .A(n6456), .B(n6794), .C(n899), .Y(n3318) );
  NAND2X1 U1676 ( .A(\Mem[32][8] ), .B(n6797), .Y(n899) );
  OAI21X1 U1677 ( .A(n6451), .B(n6794), .C(n900), .Y(n3319) );
  NAND2X1 U1678 ( .A(\Mem[32][9] ), .B(n6797), .Y(n900) );
  OAI21X1 U1679 ( .A(n6601), .B(n6794), .C(n901), .Y(n3320) );
  NAND2X1 U1680 ( .A(\Mem[32][10] ), .B(n6797), .Y(n901) );
  OAI21X1 U1681 ( .A(n6596), .B(n6794), .C(n902), .Y(n3321) );
  NAND2X1 U1682 ( .A(\Mem[32][11] ), .B(n6797), .Y(n902) );
  OAI21X1 U1683 ( .A(n6591), .B(n6794), .C(n903), .Y(n3322) );
  NAND2X1 U1684 ( .A(\Mem[32][12] ), .B(n6797), .Y(n903) );
  OAI21X1 U1685 ( .A(n6586), .B(n6795), .C(n904), .Y(n3323) );
  NAND2X1 U1686 ( .A(\Mem[32][13] ), .B(n6797), .Y(n904) );
  OAI21X1 U1687 ( .A(n6581), .B(n6795), .C(n905), .Y(n3324) );
  NAND2X1 U1688 ( .A(\Mem[32][14] ), .B(n6797), .Y(n905) );
  OAI21X1 U1689 ( .A(n6576), .B(n6795), .C(n906), .Y(n3325) );
  NAND2X1 U1690 ( .A(\Mem[32][15] ), .B(n6796), .Y(n906) );
  OAI21X1 U1691 ( .A(n6571), .B(n6795), .C(n907), .Y(n3326) );
  NAND2X1 U1692 ( .A(\Mem[32][16] ), .B(n6797), .Y(n907) );
  OAI21X1 U1693 ( .A(n6566), .B(n6795), .C(n908), .Y(n3327) );
  NAND2X1 U1694 ( .A(\Mem[32][17] ), .B(n6796), .Y(n908) );
  OAI21X1 U1695 ( .A(n6561), .B(n6795), .C(n909), .Y(n3328) );
  NAND2X1 U1696 ( .A(\Mem[32][18] ), .B(n6796), .Y(n909) );
  OAI21X1 U1697 ( .A(n6556), .B(n6795), .C(n910), .Y(n3329) );
  NAND2X1 U1698 ( .A(\Mem[32][19] ), .B(n6796), .Y(n910) );
  OAI21X1 U1699 ( .A(n6546), .B(n6795), .C(n911), .Y(n3330) );
  NAND2X1 U1700 ( .A(\Mem[32][20] ), .B(n6796), .Y(n911) );
  OAI21X1 U1701 ( .A(n6541), .B(n6795), .C(n912), .Y(n3331) );
  NAND2X1 U1702 ( .A(\Mem[32][21] ), .B(n6796), .Y(n912) );
  OAI21X1 U1703 ( .A(n6536), .B(n6795), .C(n913), .Y(n3332) );
  NAND2X1 U1704 ( .A(\Mem[32][22] ), .B(n6797), .Y(n913) );
  OAI21X1 U1705 ( .A(n6531), .B(n6796), .C(n914), .Y(n3333) );
  NAND2X1 U1706 ( .A(\Mem[32][23] ), .B(n6796), .Y(n914) );
  OAI21X1 U1707 ( .A(n6526), .B(n6795), .C(n915), .Y(n3334) );
  NAND2X1 U1708 ( .A(\Mem[32][24] ), .B(n6797), .Y(n915) );
  OAI21X1 U1709 ( .A(n6521), .B(n6796), .C(n916), .Y(n3335) );
  NAND2X1 U1710 ( .A(\Mem[32][25] ), .B(n6797), .Y(n916) );
  OAI21X1 U1711 ( .A(n6516), .B(n6796), .C(n917), .Y(n3336) );
  NAND2X1 U1712 ( .A(\Mem[32][26] ), .B(n6797), .Y(n917) );
  OAI21X1 U1713 ( .A(n6511), .B(n6796), .C(n918), .Y(n3337) );
  NAND2X1 U1714 ( .A(\Mem[32][27] ), .B(n6797), .Y(n918) );
  OAI21X1 U1715 ( .A(n6506), .B(n6796), .C(n919), .Y(n3338) );
  NAND2X1 U1716 ( .A(\Mem[32][28] ), .B(n6797), .Y(n919) );
  OAI21X1 U1717 ( .A(n6501), .B(n6796), .C(n920), .Y(n3339) );
  NAND2X1 U1718 ( .A(\Mem[32][29] ), .B(n6797), .Y(n920) );
  OAI21X1 U1719 ( .A(n6491), .B(n6796), .C(n921), .Y(n3340) );
  NAND2X1 U1720 ( .A(\Mem[32][30] ), .B(n6798), .Y(n921) );
  OAI21X1 U1721 ( .A(n6486), .B(n6796), .C(n922), .Y(n3341) );
  NAND2X1 U1722 ( .A(\Mem[32][31] ), .B(n6798), .Y(n922) );
  NAND2X1 U1723 ( .A(n7011), .B(n7016), .Y(n890) );
  OAI21X1 U1724 ( .A(n6606), .B(n6790), .C(n925), .Y(n3342) );
  NAND2X1 U1725 ( .A(\Mem[33][0] ), .B(n6793), .Y(n925) );
  OAI21X1 U1726 ( .A(n6551), .B(n6789), .C(n926), .Y(n3343) );
  NAND2X1 U1727 ( .A(\Mem[33][1] ), .B(n6793), .Y(n926) );
  OAI21X1 U1728 ( .A(n6496), .B(n6789), .C(n927), .Y(n3344) );
  NAND2X1 U1729 ( .A(\Mem[33][2] ), .B(n6793), .Y(n927) );
  OAI21X1 U1730 ( .A(n6481), .B(n6789), .C(n928), .Y(n3345) );
  NAND2X1 U1731 ( .A(\Mem[33][3] ), .B(n6792), .Y(n928) );
  OAI21X1 U1732 ( .A(n6476), .B(n6789), .C(n929), .Y(n3346) );
  NAND2X1 U1733 ( .A(\Mem[33][4] ), .B(n6793), .Y(n929) );
  OAI21X1 U1734 ( .A(n6471), .B(n6789), .C(n930), .Y(n3347) );
  NAND2X1 U1735 ( .A(\Mem[33][5] ), .B(n6792), .Y(n930) );
  OAI21X1 U1736 ( .A(n6466), .B(n6789), .C(n931), .Y(n3348) );
  NAND2X1 U1737 ( .A(\Mem[33][6] ), .B(n6792), .Y(n931) );
  OAI21X1 U1738 ( .A(n6461), .B(n6789), .C(n932), .Y(n3349) );
  NAND2X1 U1739 ( .A(\Mem[33][7] ), .B(n6792), .Y(n932) );
  OAI21X1 U1740 ( .A(n6456), .B(n6789), .C(n933), .Y(n3350) );
  NAND2X1 U1741 ( .A(\Mem[33][8] ), .B(n6792), .Y(n933) );
  OAI21X1 U1742 ( .A(n6451), .B(n6789), .C(n934), .Y(n3351) );
  NAND2X1 U1743 ( .A(\Mem[33][9] ), .B(n6792), .Y(n934) );
  OAI21X1 U1744 ( .A(n6601), .B(n6789), .C(n935), .Y(n3352) );
  NAND2X1 U1745 ( .A(\Mem[33][10] ), .B(n6792), .Y(n935) );
  OAI21X1 U1746 ( .A(n6596), .B(n6789), .C(n936), .Y(n3353) );
  NAND2X1 U1747 ( .A(\Mem[33][11] ), .B(n6792), .Y(n936) );
  OAI21X1 U1748 ( .A(n6591), .B(n6789), .C(n937), .Y(n3354) );
  NAND2X1 U1749 ( .A(\Mem[33][12] ), .B(n6792), .Y(n937) );
  OAI21X1 U1750 ( .A(n6586), .B(n6790), .C(n938), .Y(n3355) );
  NAND2X1 U1751 ( .A(\Mem[33][13] ), .B(n6792), .Y(n938) );
  OAI21X1 U1752 ( .A(n6581), .B(n6790), .C(n939), .Y(n3356) );
  NAND2X1 U1753 ( .A(\Mem[33][14] ), .B(n6792), .Y(n939) );
  OAI21X1 U1754 ( .A(n6576), .B(n6790), .C(n940), .Y(n3357) );
  NAND2X1 U1755 ( .A(\Mem[33][15] ), .B(n6791), .Y(n940) );
  OAI21X1 U1756 ( .A(n6571), .B(n6790), .C(n941), .Y(n3358) );
  NAND2X1 U1757 ( .A(\Mem[33][16] ), .B(n6792), .Y(n941) );
  OAI21X1 U1758 ( .A(n6566), .B(n6790), .C(n942), .Y(n3359) );
  NAND2X1 U1759 ( .A(\Mem[33][17] ), .B(n6791), .Y(n942) );
  OAI21X1 U1760 ( .A(n6561), .B(n6790), .C(n943), .Y(n3360) );
  NAND2X1 U1761 ( .A(\Mem[33][18] ), .B(n6791), .Y(n943) );
  OAI21X1 U1762 ( .A(n6556), .B(n6790), .C(n944), .Y(n3361) );
  NAND2X1 U1763 ( .A(\Mem[33][19] ), .B(n6791), .Y(n944) );
  OAI21X1 U1764 ( .A(n6546), .B(n6790), .C(n945), .Y(n3362) );
  NAND2X1 U1765 ( .A(\Mem[33][20] ), .B(n6791), .Y(n945) );
  OAI21X1 U1766 ( .A(n6541), .B(n6790), .C(n946), .Y(n3363) );
  NAND2X1 U1767 ( .A(\Mem[33][21] ), .B(n6791), .Y(n946) );
  OAI21X1 U1768 ( .A(n6536), .B(n6790), .C(n947), .Y(n3364) );
  NAND2X1 U1769 ( .A(\Mem[33][22] ), .B(n6792), .Y(n947) );
  OAI21X1 U1770 ( .A(n6531), .B(n6791), .C(n948), .Y(n3365) );
  NAND2X1 U1771 ( .A(\Mem[33][23] ), .B(n6791), .Y(n948) );
  OAI21X1 U1772 ( .A(n6526), .B(n6790), .C(n949), .Y(n3366) );
  NAND2X1 U1773 ( .A(\Mem[33][24] ), .B(n6792), .Y(n949) );
  OAI21X1 U1774 ( .A(n6521), .B(n6791), .C(n950), .Y(n3367) );
  NAND2X1 U1775 ( .A(\Mem[33][25] ), .B(n6792), .Y(n950) );
  OAI21X1 U1776 ( .A(n6516), .B(n6791), .C(n951), .Y(n3368) );
  NAND2X1 U1777 ( .A(\Mem[33][26] ), .B(n6792), .Y(n951) );
  OAI21X1 U1778 ( .A(n6511), .B(n6791), .C(n952), .Y(n3369) );
  NAND2X1 U1779 ( .A(\Mem[33][27] ), .B(n6792), .Y(n952) );
  OAI21X1 U1780 ( .A(n6506), .B(n6791), .C(n953), .Y(n3370) );
  NAND2X1 U1781 ( .A(\Mem[33][28] ), .B(n6792), .Y(n953) );
  OAI21X1 U1782 ( .A(n6501), .B(n6791), .C(n954), .Y(n3371) );
  NAND2X1 U1783 ( .A(\Mem[33][29] ), .B(n6792), .Y(n954) );
  OAI21X1 U1784 ( .A(n6491), .B(n6791), .C(n955), .Y(n3372) );
  NAND2X1 U1785 ( .A(\Mem[33][30] ), .B(n6793), .Y(n955) );
  OAI21X1 U1786 ( .A(n6486), .B(n6791), .C(n956), .Y(n3373) );
  NAND2X1 U1787 ( .A(\Mem[33][31] ), .B(n6793), .Y(n956) );
  NAND2X1 U1788 ( .A(n7011), .B(n7017), .Y(n924) );
  OAI21X1 U1789 ( .A(n6606), .B(n6785), .C(n958), .Y(n3374) );
  NAND2X1 U1790 ( .A(\Mem[34][0] ), .B(n6788), .Y(n958) );
  OAI21X1 U1791 ( .A(n6551), .B(n6784), .C(n959), .Y(n3375) );
  NAND2X1 U1792 ( .A(\Mem[34][1] ), .B(n6788), .Y(n959) );
  OAI21X1 U1793 ( .A(n6496), .B(n6784), .C(n960), .Y(n3376) );
  NAND2X1 U1794 ( .A(\Mem[34][2] ), .B(n6788), .Y(n960) );
  OAI21X1 U1795 ( .A(n6481), .B(n6784), .C(n961), .Y(n3377) );
  NAND2X1 U1796 ( .A(\Mem[34][3] ), .B(n6787), .Y(n961) );
  OAI21X1 U1797 ( .A(n6476), .B(n6784), .C(n962), .Y(n3378) );
  NAND2X1 U1798 ( .A(\Mem[34][4] ), .B(n6788), .Y(n962) );
  OAI21X1 U1799 ( .A(n6471), .B(n6784), .C(n963), .Y(n3379) );
  NAND2X1 U1800 ( .A(\Mem[34][5] ), .B(n6787), .Y(n963) );
  OAI21X1 U1801 ( .A(n6466), .B(n6784), .C(n964), .Y(n3380) );
  NAND2X1 U1802 ( .A(\Mem[34][6] ), .B(n6787), .Y(n964) );
  OAI21X1 U1803 ( .A(n6461), .B(n6784), .C(n965), .Y(n3381) );
  NAND2X1 U1804 ( .A(\Mem[34][7] ), .B(n6787), .Y(n965) );
  OAI21X1 U1805 ( .A(n6456), .B(n6784), .C(n966), .Y(n3382) );
  NAND2X1 U1806 ( .A(\Mem[34][8] ), .B(n6787), .Y(n966) );
  OAI21X1 U1807 ( .A(n6451), .B(n6784), .C(n967), .Y(n3383) );
  NAND2X1 U1808 ( .A(\Mem[34][9] ), .B(n6787), .Y(n967) );
  OAI21X1 U1809 ( .A(n6601), .B(n6784), .C(n968), .Y(n3384) );
  NAND2X1 U1810 ( .A(\Mem[34][10] ), .B(n6787), .Y(n968) );
  OAI21X1 U1811 ( .A(n6596), .B(n6784), .C(n969), .Y(n3385) );
  NAND2X1 U1812 ( .A(\Mem[34][11] ), .B(n6787), .Y(n969) );
  OAI21X1 U1813 ( .A(n6591), .B(n6784), .C(n970), .Y(n3386) );
  NAND2X1 U1814 ( .A(\Mem[34][12] ), .B(n6787), .Y(n970) );
  OAI21X1 U1815 ( .A(n6586), .B(n6785), .C(n971), .Y(n3387) );
  NAND2X1 U1816 ( .A(\Mem[34][13] ), .B(n6787), .Y(n971) );
  OAI21X1 U1817 ( .A(n6581), .B(n6785), .C(n972), .Y(n3388) );
  NAND2X1 U1818 ( .A(\Mem[34][14] ), .B(n6787), .Y(n972) );
  OAI21X1 U1819 ( .A(n6576), .B(n6785), .C(n973), .Y(n3389) );
  NAND2X1 U1820 ( .A(\Mem[34][15] ), .B(n6786), .Y(n973) );
  OAI21X1 U1821 ( .A(n6571), .B(n6785), .C(n974), .Y(n3390) );
  NAND2X1 U1822 ( .A(\Mem[34][16] ), .B(n6787), .Y(n974) );
  OAI21X1 U1823 ( .A(n6566), .B(n6785), .C(n975), .Y(n3391) );
  NAND2X1 U1824 ( .A(\Mem[34][17] ), .B(n6786), .Y(n975) );
  OAI21X1 U1825 ( .A(n6561), .B(n6785), .C(n976), .Y(n3392) );
  NAND2X1 U1826 ( .A(\Mem[34][18] ), .B(n6786), .Y(n976) );
  OAI21X1 U1827 ( .A(n6556), .B(n6785), .C(n977), .Y(n3393) );
  NAND2X1 U1828 ( .A(\Mem[34][19] ), .B(n6786), .Y(n977) );
  OAI21X1 U1829 ( .A(n6546), .B(n6785), .C(n978), .Y(n3394) );
  NAND2X1 U1830 ( .A(\Mem[34][20] ), .B(n6786), .Y(n978) );
  OAI21X1 U1831 ( .A(n6541), .B(n6785), .C(n979), .Y(n3395) );
  NAND2X1 U1832 ( .A(\Mem[34][21] ), .B(n6786), .Y(n979) );
  OAI21X1 U1833 ( .A(n6536), .B(n6785), .C(n980), .Y(n3396) );
  NAND2X1 U1834 ( .A(\Mem[34][22] ), .B(n6787), .Y(n980) );
  OAI21X1 U1835 ( .A(n6531), .B(n6786), .C(n981), .Y(n3397) );
  NAND2X1 U1836 ( .A(\Mem[34][23] ), .B(n6786), .Y(n981) );
  OAI21X1 U1837 ( .A(n6526), .B(n6785), .C(n982), .Y(n3398) );
  NAND2X1 U1838 ( .A(\Mem[34][24] ), .B(n6787), .Y(n982) );
  OAI21X1 U1839 ( .A(n6521), .B(n6786), .C(n983), .Y(n3399) );
  NAND2X1 U1840 ( .A(\Mem[34][25] ), .B(n6787), .Y(n983) );
  OAI21X1 U1841 ( .A(n6516), .B(n6786), .C(n984), .Y(n3400) );
  NAND2X1 U1842 ( .A(\Mem[34][26] ), .B(n6787), .Y(n984) );
  OAI21X1 U1843 ( .A(n6511), .B(n6786), .C(n985), .Y(n3401) );
  NAND2X1 U1844 ( .A(\Mem[34][27] ), .B(n6787), .Y(n985) );
  OAI21X1 U1845 ( .A(n6506), .B(n6786), .C(n986), .Y(n3402) );
  NAND2X1 U1846 ( .A(\Mem[34][28] ), .B(n6787), .Y(n986) );
  OAI21X1 U1847 ( .A(n6501), .B(n6786), .C(n987), .Y(n3403) );
  NAND2X1 U1848 ( .A(\Mem[34][29] ), .B(n6787), .Y(n987) );
  OAI21X1 U1849 ( .A(n6491), .B(n6786), .C(n988), .Y(n3404) );
  NAND2X1 U1850 ( .A(\Mem[34][30] ), .B(n6788), .Y(n988) );
  OAI21X1 U1851 ( .A(n6486), .B(n6786), .C(n989), .Y(n3405) );
  NAND2X1 U1852 ( .A(\Mem[34][31] ), .B(n6788), .Y(n989) );
  NAND2X1 U1853 ( .A(n7011), .B(n7018), .Y(n957) );
  OAI21X1 U1854 ( .A(n6606), .B(n6780), .C(n991), .Y(n3406) );
  NAND2X1 U1855 ( .A(\Mem[35][0] ), .B(n6783), .Y(n991) );
  OAI21X1 U1856 ( .A(n6551), .B(n6779), .C(n992), .Y(n3407) );
  NAND2X1 U1857 ( .A(\Mem[35][1] ), .B(n6783), .Y(n992) );
  OAI21X1 U1858 ( .A(n6496), .B(n6779), .C(n993), .Y(n3408) );
  NAND2X1 U1859 ( .A(\Mem[35][2] ), .B(n6783), .Y(n993) );
  OAI21X1 U1860 ( .A(n6481), .B(n6779), .C(n994), .Y(n3409) );
  NAND2X1 U1861 ( .A(\Mem[35][3] ), .B(n6782), .Y(n994) );
  OAI21X1 U1862 ( .A(n6476), .B(n6779), .C(n995), .Y(n3410) );
  NAND2X1 U1863 ( .A(\Mem[35][4] ), .B(n6783), .Y(n995) );
  OAI21X1 U1864 ( .A(n6471), .B(n6779), .C(n996), .Y(n3411) );
  NAND2X1 U1865 ( .A(\Mem[35][5] ), .B(n6782), .Y(n996) );
  OAI21X1 U1866 ( .A(n6466), .B(n6779), .C(n997), .Y(n3412) );
  NAND2X1 U1867 ( .A(\Mem[35][6] ), .B(n6782), .Y(n997) );
  OAI21X1 U1868 ( .A(n6461), .B(n6779), .C(n998), .Y(n3413) );
  NAND2X1 U1869 ( .A(\Mem[35][7] ), .B(n6782), .Y(n998) );
  OAI21X1 U1870 ( .A(n6456), .B(n6779), .C(n999), .Y(n3414) );
  NAND2X1 U1871 ( .A(\Mem[35][8] ), .B(n6782), .Y(n999) );
  OAI21X1 U1872 ( .A(n6451), .B(n6779), .C(n1000), .Y(n3415) );
  NAND2X1 U1873 ( .A(\Mem[35][9] ), .B(n6782), .Y(n1000) );
  OAI21X1 U1874 ( .A(n6601), .B(n6779), .C(n1001), .Y(n3416) );
  NAND2X1 U1875 ( .A(\Mem[35][10] ), .B(n6782), .Y(n1001) );
  OAI21X1 U1876 ( .A(n6596), .B(n6779), .C(n1002), .Y(n3417) );
  NAND2X1 U1877 ( .A(\Mem[35][11] ), .B(n6782), .Y(n1002) );
  OAI21X1 U1878 ( .A(n6591), .B(n6779), .C(n1003), .Y(n3418) );
  NAND2X1 U1879 ( .A(\Mem[35][12] ), .B(n6782), .Y(n1003) );
  OAI21X1 U1880 ( .A(n6586), .B(n6780), .C(n1004), .Y(n3419) );
  NAND2X1 U1881 ( .A(\Mem[35][13] ), .B(n6782), .Y(n1004) );
  OAI21X1 U1882 ( .A(n6581), .B(n6780), .C(n1005), .Y(n3420) );
  NAND2X1 U1883 ( .A(\Mem[35][14] ), .B(n6782), .Y(n1005) );
  OAI21X1 U1884 ( .A(n6576), .B(n6780), .C(n1006), .Y(n3421) );
  NAND2X1 U1885 ( .A(\Mem[35][15] ), .B(n6781), .Y(n1006) );
  OAI21X1 U1886 ( .A(n6571), .B(n6780), .C(n1007), .Y(n3422) );
  NAND2X1 U1887 ( .A(\Mem[35][16] ), .B(n6782), .Y(n1007) );
  OAI21X1 U1888 ( .A(n6566), .B(n6780), .C(n1008), .Y(n3423) );
  NAND2X1 U1889 ( .A(\Mem[35][17] ), .B(n6781), .Y(n1008) );
  OAI21X1 U1890 ( .A(n6561), .B(n6780), .C(n1009), .Y(n3424) );
  NAND2X1 U1891 ( .A(\Mem[35][18] ), .B(n6781), .Y(n1009) );
  OAI21X1 U1892 ( .A(n6556), .B(n6780), .C(n1010), .Y(n3425) );
  NAND2X1 U1893 ( .A(\Mem[35][19] ), .B(n6781), .Y(n1010) );
  OAI21X1 U1894 ( .A(n6546), .B(n6780), .C(n1011), .Y(n3426) );
  NAND2X1 U1895 ( .A(\Mem[35][20] ), .B(n6781), .Y(n1011) );
  OAI21X1 U1896 ( .A(n6541), .B(n6780), .C(n1012), .Y(n3427) );
  NAND2X1 U1897 ( .A(\Mem[35][21] ), .B(n6781), .Y(n1012) );
  OAI21X1 U1898 ( .A(n6536), .B(n6780), .C(n1013), .Y(n3428) );
  NAND2X1 U1899 ( .A(\Mem[35][22] ), .B(n6782), .Y(n1013) );
  OAI21X1 U1900 ( .A(n6531), .B(n6781), .C(n1014), .Y(n3429) );
  NAND2X1 U1901 ( .A(\Mem[35][23] ), .B(n6781), .Y(n1014) );
  OAI21X1 U1902 ( .A(n6526), .B(n6780), .C(n1015), .Y(n3430) );
  NAND2X1 U1903 ( .A(\Mem[35][24] ), .B(n6782), .Y(n1015) );
  OAI21X1 U1904 ( .A(n6521), .B(n6781), .C(n1016), .Y(n3431) );
  NAND2X1 U1905 ( .A(\Mem[35][25] ), .B(n6782), .Y(n1016) );
  OAI21X1 U1906 ( .A(n6516), .B(n6781), .C(n1017), .Y(n3432) );
  NAND2X1 U1907 ( .A(\Mem[35][26] ), .B(n6782), .Y(n1017) );
  OAI21X1 U1908 ( .A(n6511), .B(n6781), .C(n1018), .Y(n3433) );
  NAND2X1 U1909 ( .A(\Mem[35][27] ), .B(n6782), .Y(n1018) );
  OAI21X1 U1910 ( .A(n6506), .B(n6781), .C(n1019), .Y(n3434) );
  NAND2X1 U1911 ( .A(\Mem[35][28] ), .B(n6782), .Y(n1019) );
  OAI21X1 U1912 ( .A(n6501), .B(n6781), .C(n1020), .Y(n3435) );
  NAND2X1 U1913 ( .A(\Mem[35][29] ), .B(n6782), .Y(n1020) );
  OAI21X1 U1914 ( .A(n6491), .B(n6781), .C(n1021), .Y(n3436) );
  NAND2X1 U1915 ( .A(\Mem[35][30] ), .B(n6783), .Y(n1021) );
  OAI21X1 U1916 ( .A(n6486), .B(n6781), .C(n1022), .Y(n3437) );
  NAND2X1 U1917 ( .A(\Mem[35][31] ), .B(n6783), .Y(n1022) );
  NAND2X1 U1918 ( .A(n7011), .B(n7019), .Y(n990) );
  OAI21X1 U1919 ( .A(n6606), .B(n6775), .C(n1024), .Y(n3438) );
  NAND2X1 U1920 ( .A(\Mem[36][0] ), .B(n6778), .Y(n1024) );
  OAI21X1 U1921 ( .A(n6551), .B(n6774), .C(n1025), .Y(n3439) );
  NAND2X1 U1922 ( .A(\Mem[36][1] ), .B(n6778), .Y(n1025) );
  OAI21X1 U1923 ( .A(n6496), .B(n6774), .C(n1026), .Y(n3440) );
  NAND2X1 U1924 ( .A(\Mem[36][2] ), .B(n6778), .Y(n1026) );
  OAI21X1 U1925 ( .A(n6481), .B(n6774), .C(n1027), .Y(n3441) );
  NAND2X1 U1926 ( .A(\Mem[36][3] ), .B(n6777), .Y(n1027) );
  OAI21X1 U1927 ( .A(n6476), .B(n6774), .C(n1028), .Y(n3442) );
  NAND2X1 U1928 ( .A(\Mem[36][4] ), .B(n6778), .Y(n1028) );
  OAI21X1 U1929 ( .A(n6471), .B(n6774), .C(n1029), .Y(n3443) );
  NAND2X1 U1930 ( .A(\Mem[36][5] ), .B(n6777), .Y(n1029) );
  OAI21X1 U1931 ( .A(n6466), .B(n6774), .C(n1030), .Y(n3444) );
  NAND2X1 U1932 ( .A(\Mem[36][6] ), .B(n6777), .Y(n1030) );
  OAI21X1 U1933 ( .A(n6461), .B(n6774), .C(n1031), .Y(n3445) );
  NAND2X1 U1934 ( .A(\Mem[36][7] ), .B(n6777), .Y(n1031) );
  OAI21X1 U1935 ( .A(n6456), .B(n6774), .C(n1032), .Y(n3446) );
  NAND2X1 U1936 ( .A(\Mem[36][8] ), .B(n6777), .Y(n1032) );
  OAI21X1 U1937 ( .A(n6451), .B(n6774), .C(n1033), .Y(n3447) );
  NAND2X1 U1938 ( .A(\Mem[36][9] ), .B(n6777), .Y(n1033) );
  OAI21X1 U1939 ( .A(n6601), .B(n6774), .C(n1034), .Y(n3448) );
  NAND2X1 U1940 ( .A(\Mem[36][10] ), .B(n6777), .Y(n1034) );
  OAI21X1 U1941 ( .A(n6596), .B(n6774), .C(n1035), .Y(n3449) );
  NAND2X1 U1942 ( .A(\Mem[36][11] ), .B(n6777), .Y(n1035) );
  OAI21X1 U1943 ( .A(n6591), .B(n6774), .C(n1036), .Y(n3450) );
  NAND2X1 U1944 ( .A(\Mem[36][12] ), .B(n6777), .Y(n1036) );
  OAI21X1 U1945 ( .A(n6586), .B(n6775), .C(n1037), .Y(n3451) );
  NAND2X1 U1946 ( .A(\Mem[36][13] ), .B(n6777), .Y(n1037) );
  OAI21X1 U1947 ( .A(n6581), .B(n6775), .C(n1038), .Y(n3452) );
  NAND2X1 U1948 ( .A(\Mem[36][14] ), .B(n6777), .Y(n1038) );
  OAI21X1 U1949 ( .A(n6576), .B(n6775), .C(n1039), .Y(n3453) );
  NAND2X1 U1950 ( .A(\Mem[36][15] ), .B(n6776), .Y(n1039) );
  OAI21X1 U1951 ( .A(n6571), .B(n6775), .C(n1040), .Y(n3454) );
  NAND2X1 U1952 ( .A(\Mem[36][16] ), .B(n6777), .Y(n1040) );
  OAI21X1 U1953 ( .A(n6566), .B(n6775), .C(n1041), .Y(n3455) );
  NAND2X1 U1954 ( .A(\Mem[36][17] ), .B(n6776), .Y(n1041) );
  OAI21X1 U1955 ( .A(n6561), .B(n6775), .C(n1042), .Y(n3456) );
  NAND2X1 U1956 ( .A(\Mem[36][18] ), .B(n6776), .Y(n1042) );
  OAI21X1 U1957 ( .A(n6556), .B(n6775), .C(n1043), .Y(n3457) );
  NAND2X1 U1958 ( .A(\Mem[36][19] ), .B(n6776), .Y(n1043) );
  OAI21X1 U1959 ( .A(n6546), .B(n6775), .C(n1044), .Y(n3458) );
  NAND2X1 U1960 ( .A(\Mem[36][20] ), .B(n6776), .Y(n1044) );
  OAI21X1 U1961 ( .A(n6541), .B(n6775), .C(n1045), .Y(n3459) );
  NAND2X1 U1962 ( .A(\Mem[36][21] ), .B(n6776), .Y(n1045) );
  OAI21X1 U1963 ( .A(n6536), .B(n6775), .C(n1046), .Y(n3460) );
  NAND2X1 U1964 ( .A(\Mem[36][22] ), .B(n6777), .Y(n1046) );
  OAI21X1 U1965 ( .A(n6531), .B(n6776), .C(n1047), .Y(n3461) );
  NAND2X1 U1966 ( .A(\Mem[36][23] ), .B(n6776), .Y(n1047) );
  OAI21X1 U1967 ( .A(n6526), .B(n6775), .C(n1048), .Y(n3462) );
  NAND2X1 U1968 ( .A(\Mem[36][24] ), .B(n6777), .Y(n1048) );
  OAI21X1 U1969 ( .A(n6521), .B(n6776), .C(n1049), .Y(n3463) );
  NAND2X1 U1970 ( .A(\Mem[36][25] ), .B(n6777), .Y(n1049) );
  OAI21X1 U1971 ( .A(n6516), .B(n6776), .C(n1050), .Y(n3464) );
  NAND2X1 U1972 ( .A(\Mem[36][26] ), .B(n6777), .Y(n1050) );
  OAI21X1 U1973 ( .A(n6511), .B(n6776), .C(n1051), .Y(n3465) );
  NAND2X1 U1974 ( .A(\Mem[36][27] ), .B(n6777), .Y(n1051) );
  OAI21X1 U1975 ( .A(n6506), .B(n6776), .C(n1052), .Y(n3466) );
  NAND2X1 U1976 ( .A(\Mem[36][28] ), .B(n6777), .Y(n1052) );
  OAI21X1 U1977 ( .A(n6501), .B(n6776), .C(n1053), .Y(n3467) );
  NAND2X1 U1978 ( .A(\Mem[36][29] ), .B(n6777), .Y(n1053) );
  OAI21X1 U1979 ( .A(n6491), .B(n6776), .C(n1054), .Y(n3468) );
  NAND2X1 U1980 ( .A(\Mem[36][30] ), .B(n6778), .Y(n1054) );
  OAI21X1 U1981 ( .A(n6486), .B(n6776), .C(n1055), .Y(n3469) );
  NAND2X1 U1982 ( .A(\Mem[36][31] ), .B(n6778), .Y(n1055) );
  NAND2X1 U1983 ( .A(n7011), .B(n7022), .Y(n1023) );
  OAI21X1 U1984 ( .A(n6606), .B(n6770), .C(n1057), .Y(n3470) );
  NAND2X1 U1985 ( .A(\Mem[37][0] ), .B(n6773), .Y(n1057) );
  OAI21X1 U1986 ( .A(n6551), .B(n6769), .C(n1058), .Y(n3471) );
  NAND2X1 U1987 ( .A(\Mem[37][1] ), .B(n6773), .Y(n1058) );
  OAI21X1 U1988 ( .A(n6496), .B(n6769), .C(n1059), .Y(n3472) );
  NAND2X1 U1989 ( .A(\Mem[37][2] ), .B(n6773), .Y(n1059) );
  OAI21X1 U1990 ( .A(n6481), .B(n6769), .C(n1060), .Y(n3473) );
  NAND2X1 U1991 ( .A(\Mem[37][3] ), .B(n6772), .Y(n1060) );
  OAI21X1 U1992 ( .A(n6476), .B(n6769), .C(n1061), .Y(n3474) );
  NAND2X1 U1993 ( .A(\Mem[37][4] ), .B(n6773), .Y(n1061) );
  OAI21X1 U1994 ( .A(n6471), .B(n6769), .C(n1062), .Y(n3475) );
  NAND2X1 U1995 ( .A(\Mem[37][5] ), .B(n6772), .Y(n1062) );
  OAI21X1 U1996 ( .A(n6466), .B(n6769), .C(n1063), .Y(n3476) );
  NAND2X1 U1997 ( .A(\Mem[37][6] ), .B(n6772), .Y(n1063) );
  OAI21X1 U1998 ( .A(n6461), .B(n6769), .C(n1064), .Y(n3477) );
  NAND2X1 U1999 ( .A(\Mem[37][7] ), .B(n6772), .Y(n1064) );
  OAI21X1 U2000 ( .A(n6456), .B(n6769), .C(n1065), .Y(n3478) );
  NAND2X1 U2001 ( .A(\Mem[37][8] ), .B(n6772), .Y(n1065) );
  OAI21X1 U2002 ( .A(n6451), .B(n6769), .C(n1066), .Y(n3479) );
  NAND2X1 U2003 ( .A(\Mem[37][9] ), .B(n6772), .Y(n1066) );
  OAI21X1 U2004 ( .A(n6601), .B(n6769), .C(n1067), .Y(n3480) );
  NAND2X1 U2005 ( .A(\Mem[37][10] ), .B(n6772), .Y(n1067) );
  OAI21X1 U2006 ( .A(n6596), .B(n6769), .C(n1068), .Y(n3481) );
  NAND2X1 U2007 ( .A(\Mem[37][11] ), .B(n6772), .Y(n1068) );
  OAI21X1 U2008 ( .A(n6591), .B(n6769), .C(n1069), .Y(n3482) );
  NAND2X1 U2009 ( .A(\Mem[37][12] ), .B(n6772), .Y(n1069) );
  OAI21X1 U2010 ( .A(n6586), .B(n6770), .C(n1070), .Y(n3483) );
  NAND2X1 U2011 ( .A(\Mem[37][13] ), .B(n6772), .Y(n1070) );
  OAI21X1 U2012 ( .A(n6581), .B(n6770), .C(n1071), .Y(n3484) );
  NAND2X1 U2013 ( .A(\Mem[37][14] ), .B(n6772), .Y(n1071) );
  OAI21X1 U2014 ( .A(n6576), .B(n6770), .C(n1072), .Y(n3485) );
  NAND2X1 U2015 ( .A(\Mem[37][15] ), .B(n6771), .Y(n1072) );
  OAI21X1 U2016 ( .A(n6571), .B(n6770), .C(n1073), .Y(n3486) );
  NAND2X1 U2017 ( .A(\Mem[37][16] ), .B(n6772), .Y(n1073) );
  OAI21X1 U2018 ( .A(n6566), .B(n6770), .C(n1074), .Y(n3487) );
  NAND2X1 U2019 ( .A(\Mem[37][17] ), .B(n6771), .Y(n1074) );
  OAI21X1 U2020 ( .A(n6561), .B(n6770), .C(n1075), .Y(n3488) );
  NAND2X1 U2021 ( .A(\Mem[37][18] ), .B(n6771), .Y(n1075) );
  OAI21X1 U2022 ( .A(n6556), .B(n6770), .C(n1076), .Y(n3489) );
  NAND2X1 U2023 ( .A(\Mem[37][19] ), .B(n6771), .Y(n1076) );
  OAI21X1 U2024 ( .A(n6546), .B(n6770), .C(n1077), .Y(n3490) );
  NAND2X1 U2025 ( .A(\Mem[37][20] ), .B(n6771), .Y(n1077) );
  OAI21X1 U2026 ( .A(n6541), .B(n6770), .C(n1078), .Y(n3491) );
  NAND2X1 U2027 ( .A(\Mem[37][21] ), .B(n6771), .Y(n1078) );
  OAI21X1 U2028 ( .A(n6536), .B(n6770), .C(n1079), .Y(n3492) );
  NAND2X1 U2029 ( .A(\Mem[37][22] ), .B(n6772), .Y(n1079) );
  OAI21X1 U2030 ( .A(n6531), .B(n6771), .C(n1080), .Y(n3493) );
  NAND2X1 U2031 ( .A(\Mem[37][23] ), .B(n6771), .Y(n1080) );
  OAI21X1 U2032 ( .A(n6526), .B(n6770), .C(n1081), .Y(n3494) );
  NAND2X1 U2033 ( .A(\Mem[37][24] ), .B(n6772), .Y(n1081) );
  OAI21X1 U2034 ( .A(n6521), .B(n6771), .C(n1082), .Y(n3495) );
  NAND2X1 U2035 ( .A(\Mem[37][25] ), .B(n6772), .Y(n1082) );
  OAI21X1 U2036 ( .A(n6516), .B(n6771), .C(n1083), .Y(n3496) );
  NAND2X1 U2037 ( .A(\Mem[37][26] ), .B(n6772), .Y(n1083) );
  OAI21X1 U2038 ( .A(n6511), .B(n6771), .C(n1084), .Y(n3497) );
  NAND2X1 U2039 ( .A(\Mem[37][27] ), .B(n6772), .Y(n1084) );
  OAI21X1 U2040 ( .A(n6506), .B(n6771), .C(n1085), .Y(n3498) );
  NAND2X1 U2041 ( .A(\Mem[37][28] ), .B(n6772), .Y(n1085) );
  OAI21X1 U2042 ( .A(n6501), .B(n6771), .C(n1086), .Y(n3499) );
  NAND2X1 U2043 ( .A(\Mem[37][29] ), .B(n6772), .Y(n1086) );
  OAI21X1 U2044 ( .A(n6491), .B(n6771), .C(n1087), .Y(n3500) );
  NAND2X1 U2045 ( .A(\Mem[37][30] ), .B(n6773), .Y(n1087) );
  OAI21X1 U2046 ( .A(n6486), .B(n6771), .C(n1088), .Y(n3501) );
  NAND2X1 U2047 ( .A(\Mem[37][31] ), .B(n6773), .Y(n1088) );
  NAND2X1 U2048 ( .A(n7011), .B(n7023), .Y(n1056) );
  OAI21X1 U2049 ( .A(n6606), .B(n6765), .C(n1090), .Y(n3502) );
  NAND2X1 U2050 ( .A(\Mem[38][0] ), .B(n6768), .Y(n1090) );
  OAI21X1 U2051 ( .A(n6551), .B(n6764), .C(n1091), .Y(n3503) );
  NAND2X1 U2052 ( .A(\Mem[38][1] ), .B(n6768), .Y(n1091) );
  OAI21X1 U2053 ( .A(n6496), .B(n6764), .C(n1092), .Y(n3504) );
  NAND2X1 U2054 ( .A(\Mem[38][2] ), .B(n6768), .Y(n1092) );
  OAI21X1 U2055 ( .A(n6481), .B(n6764), .C(n1093), .Y(n3505) );
  NAND2X1 U2056 ( .A(\Mem[38][3] ), .B(n6767), .Y(n1093) );
  OAI21X1 U2057 ( .A(n6476), .B(n6764), .C(n1094), .Y(n3506) );
  NAND2X1 U2058 ( .A(\Mem[38][4] ), .B(n6768), .Y(n1094) );
  OAI21X1 U2059 ( .A(n6471), .B(n6764), .C(n1095), .Y(n3507) );
  NAND2X1 U2060 ( .A(\Mem[38][5] ), .B(n6767), .Y(n1095) );
  OAI21X1 U2061 ( .A(n6466), .B(n6764), .C(n1096), .Y(n3508) );
  NAND2X1 U2062 ( .A(\Mem[38][6] ), .B(n6767), .Y(n1096) );
  OAI21X1 U2063 ( .A(n6461), .B(n6764), .C(n1097), .Y(n3509) );
  NAND2X1 U2064 ( .A(\Mem[38][7] ), .B(n6767), .Y(n1097) );
  OAI21X1 U2065 ( .A(n6456), .B(n6764), .C(n1098), .Y(n3510) );
  NAND2X1 U2066 ( .A(\Mem[38][8] ), .B(n6767), .Y(n1098) );
  OAI21X1 U2067 ( .A(n6451), .B(n6764), .C(n1099), .Y(n3511) );
  NAND2X1 U2068 ( .A(\Mem[38][9] ), .B(n6767), .Y(n1099) );
  OAI21X1 U2069 ( .A(n6601), .B(n6764), .C(n1100), .Y(n3512) );
  NAND2X1 U2070 ( .A(\Mem[38][10] ), .B(n6767), .Y(n1100) );
  OAI21X1 U2071 ( .A(n6596), .B(n6764), .C(n1101), .Y(n3513) );
  NAND2X1 U2072 ( .A(\Mem[38][11] ), .B(n6767), .Y(n1101) );
  OAI21X1 U2073 ( .A(n6591), .B(n6764), .C(n1102), .Y(n3514) );
  NAND2X1 U2074 ( .A(\Mem[38][12] ), .B(n6767), .Y(n1102) );
  OAI21X1 U2075 ( .A(n6586), .B(n6765), .C(n1103), .Y(n3515) );
  NAND2X1 U2076 ( .A(\Mem[38][13] ), .B(n6767), .Y(n1103) );
  OAI21X1 U2077 ( .A(n6581), .B(n6765), .C(n1104), .Y(n3516) );
  NAND2X1 U2078 ( .A(\Mem[38][14] ), .B(n6767), .Y(n1104) );
  OAI21X1 U2079 ( .A(n6576), .B(n6765), .C(n1105), .Y(n3517) );
  NAND2X1 U2080 ( .A(\Mem[38][15] ), .B(n6766), .Y(n1105) );
  OAI21X1 U2081 ( .A(n6571), .B(n6765), .C(n1106), .Y(n3518) );
  NAND2X1 U2082 ( .A(\Mem[38][16] ), .B(n6767), .Y(n1106) );
  OAI21X1 U2083 ( .A(n6566), .B(n6765), .C(n1107), .Y(n3519) );
  NAND2X1 U2084 ( .A(\Mem[38][17] ), .B(n6766), .Y(n1107) );
  OAI21X1 U2085 ( .A(n6561), .B(n6765), .C(n1108), .Y(n3520) );
  NAND2X1 U2086 ( .A(\Mem[38][18] ), .B(n6766), .Y(n1108) );
  OAI21X1 U2087 ( .A(n6556), .B(n6765), .C(n1109), .Y(n3521) );
  NAND2X1 U2088 ( .A(\Mem[38][19] ), .B(n6766), .Y(n1109) );
  OAI21X1 U2089 ( .A(n6546), .B(n6765), .C(n1110), .Y(n3522) );
  NAND2X1 U2090 ( .A(\Mem[38][20] ), .B(n6766), .Y(n1110) );
  OAI21X1 U2091 ( .A(n6541), .B(n6765), .C(n1111), .Y(n3523) );
  NAND2X1 U2092 ( .A(\Mem[38][21] ), .B(n6766), .Y(n1111) );
  OAI21X1 U2093 ( .A(n6536), .B(n6765), .C(n1112), .Y(n3524) );
  NAND2X1 U2094 ( .A(\Mem[38][22] ), .B(n6767), .Y(n1112) );
  OAI21X1 U2095 ( .A(n6531), .B(n6766), .C(n1113), .Y(n3525) );
  NAND2X1 U2096 ( .A(\Mem[38][23] ), .B(n6766), .Y(n1113) );
  OAI21X1 U2097 ( .A(n6526), .B(n6765), .C(n1114), .Y(n3526) );
  NAND2X1 U2098 ( .A(\Mem[38][24] ), .B(n6767), .Y(n1114) );
  OAI21X1 U2099 ( .A(n6521), .B(n6766), .C(n1115), .Y(n3527) );
  NAND2X1 U2100 ( .A(\Mem[38][25] ), .B(n6767), .Y(n1115) );
  OAI21X1 U2101 ( .A(n6516), .B(n6766), .C(n1116), .Y(n3528) );
  NAND2X1 U2102 ( .A(\Mem[38][26] ), .B(n6767), .Y(n1116) );
  OAI21X1 U2103 ( .A(n6511), .B(n6766), .C(n1117), .Y(n3529) );
  NAND2X1 U2104 ( .A(\Mem[38][27] ), .B(n6767), .Y(n1117) );
  OAI21X1 U2105 ( .A(n6506), .B(n6766), .C(n1118), .Y(n3530) );
  NAND2X1 U2106 ( .A(\Mem[38][28] ), .B(n6767), .Y(n1118) );
  OAI21X1 U2107 ( .A(n6501), .B(n6766), .C(n1119), .Y(n3531) );
  NAND2X1 U2108 ( .A(\Mem[38][29] ), .B(n6767), .Y(n1119) );
  OAI21X1 U2109 ( .A(n6491), .B(n6766), .C(n1120), .Y(n3532) );
  NAND2X1 U2110 ( .A(\Mem[38][30] ), .B(n6768), .Y(n1120) );
  OAI21X1 U2111 ( .A(n6486), .B(n6766), .C(n1121), .Y(n3533) );
  NAND2X1 U2112 ( .A(\Mem[38][31] ), .B(n6768), .Y(n1121) );
  NAND2X1 U2113 ( .A(n7011), .B(n7024), .Y(n1089) );
  OAI21X1 U2114 ( .A(n6606), .B(n6760), .C(n1123), .Y(n3534) );
  NAND2X1 U2115 ( .A(\Mem[39][0] ), .B(n6763), .Y(n1123) );
  OAI21X1 U2116 ( .A(n6551), .B(n6759), .C(n1124), .Y(n3535) );
  NAND2X1 U2117 ( .A(\Mem[39][1] ), .B(n6763), .Y(n1124) );
  OAI21X1 U2118 ( .A(n6496), .B(n6759), .C(n1125), .Y(n3536) );
  NAND2X1 U2119 ( .A(\Mem[39][2] ), .B(n6763), .Y(n1125) );
  OAI21X1 U2120 ( .A(n6481), .B(n6759), .C(n1126), .Y(n3537) );
  NAND2X1 U2121 ( .A(\Mem[39][3] ), .B(n6762), .Y(n1126) );
  OAI21X1 U2122 ( .A(n6476), .B(n6759), .C(n1127), .Y(n3538) );
  NAND2X1 U2123 ( .A(\Mem[39][4] ), .B(n6763), .Y(n1127) );
  OAI21X1 U2124 ( .A(n6471), .B(n6759), .C(n1128), .Y(n3539) );
  NAND2X1 U2125 ( .A(\Mem[39][5] ), .B(n6762), .Y(n1128) );
  OAI21X1 U2126 ( .A(n6466), .B(n6759), .C(n1129), .Y(n3540) );
  NAND2X1 U2127 ( .A(\Mem[39][6] ), .B(n6762), .Y(n1129) );
  OAI21X1 U2128 ( .A(n6461), .B(n6759), .C(n1130), .Y(n3541) );
  NAND2X1 U2129 ( .A(\Mem[39][7] ), .B(n6762), .Y(n1130) );
  OAI21X1 U2130 ( .A(n6456), .B(n6759), .C(n1131), .Y(n3542) );
  NAND2X1 U2131 ( .A(\Mem[39][8] ), .B(n6762), .Y(n1131) );
  OAI21X1 U2132 ( .A(n6451), .B(n6759), .C(n1132), .Y(n3543) );
  NAND2X1 U2133 ( .A(\Mem[39][9] ), .B(n6762), .Y(n1132) );
  OAI21X1 U2134 ( .A(n6601), .B(n6759), .C(n1133), .Y(n3544) );
  NAND2X1 U2135 ( .A(\Mem[39][10] ), .B(n6762), .Y(n1133) );
  OAI21X1 U2136 ( .A(n6596), .B(n6759), .C(n1134), .Y(n3545) );
  NAND2X1 U2137 ( .A(\Mem[39][11] ), .B(n6762), .Y(n1134) );
  OAI21X1 U2138 ( .A(n6591), .B(n6759), .C(n1135), .Y(n3546) );
  NAND2X1 U2139 ( .A(\Mem[39][12] ), .B(n6762), .Y(n1135) );
  OAI21X1 U2140 ( .A(n6586), .B(n6760), .C(n1136), .Y(n3547) );
  NAND2X1 U2141 ( .A(\Mem[39][13] ), .B(n6762), .Y(n1136) );
  OAI21X1 U2142 ( .A(n6581), .B(n6760), .C(n1137), .Y(n3548) );
  NAND2X1 U2143 ( .A(\Mem[39][14] ), .B(n6762), .Y(n1137) );
  OAI21X1 U2144 ( .A(n6576), .B(n6760), .C(n1138), .Y(n3549) );
  NAND2X1 U2145 ( .A(\Mem[39][15] ), .B(n6761), .Y(n1138) );
  OAI21X1 U2146 ( .A(n6571), .B(n6760), .C(n1139), .Y(n3550) );
  NAND2X1 U2147 ( .A(\Mem[39][16] ), .B(n6762), .Y(n1139) );
  OAI21X1 U2148 ( .A(n6566), .B(n6760), .C(n1140), .Y(n3551) );
  NAND2X1 U2149 ( .A(\Mem[39][17] ), .B(n6761), .Y(n1140) );
  OAI21X1 U2150 ( .A(n6561), .B(n6760), .C(n1141), .Y(n3552) );
  NAND2X1 U2151 ( .A(\Mem[39][18] ), .B(n6761), .Y(n1141) );
  OAI21X1 U2152 ( .A(n6556), .B(n6760), .C(n1142), .Y(n3553) );
  NAND2X1 U2153 ( .A(\Mem[39][19] ), .B(n6761), .Y(n1142) );
  OAI21X1 U2154 ( .A(n6546), .B(n6760), .C(n1143), .Y(n3554) );
  NAND2X1 U2155 ( .A(\Mem[39][20] ), .B(n6761), .Y(n1143) );
  OAI21X1 U2156 ( .A(n6541), .B(n6760), .C(n1144), .Y(n3555) );
  NAND2X1 U2157 ( .A(\Mem[39][21] ), .B(n6761), .Y(n1144) );
  OAI21X1 U2158 ( .A(n6536), .B(n6760), .C(n1145), .Y(n3556) );
  NAND2X1 U2159 ( .A(\Mem[39][22] ), .B(n6762), .Y(n1145) );
  OAI21X1 U2160 ( .A(n6531), .B(n6761), .C(n1146), .Y(n3557) );
  NAND2X1 U2161 ( .A(\Mem[39][23] ), .B(n6761), .Y(n1146) );
  OAI21X1 U2162 ( .A(n6526), .B(n6760), .C(n1147), .Y(n3558) );
  NAND2X1 U2163 ( .A(\Mem[39][24] ), .B(n6762), .Y(n1147) );
  OAI21X1 U2164 ( .A(n6521), .B(n6761), .C(n1148), .Y(n3559) );
  NAND2X1 U2165 ( .A(\Mem[39][25] ), .B(n6762), .Y(n1148) );
  OAI21X1 U2166 ( .A(n6516), .B(n6761), .C(n1149), .Y(n3560) );
  NAND2X1 U2167 ( .A(\Mem[39][26] ), .B(n6762), .Y(n1149) );
  OAI21X1 U2168 ( .A(n6511), .B(n6761), .C(n1150), .Y(n3561) );
  NAND2X1 U2169 ( .A(\Mem[39][27] ), .B(n6762), .Y(n1150) );
  OAI21X1 U2170 ( .A(n6506), .B(n6761), .C(n1151), .Y(n3562) );
  NAND2X1 U2171 ( .A(\Mem[39][28] ), .B(n6762), .Y(n1151) );
  OAI21X1 U2172 ( .A(n6501), .B(n6761), .C(n1152), .Y(n3563) );
  NAND2X1 U2173 ( .A(\Mem[39][29] ), .B(n6762), .Y(n1152) );
  OAI21X1 U2174 ( .A(n6491), .B(n6761), .C(n1153), .Y(n3564) );
  NAND2X1 U2175 ( .A(\Mem[39][30] ), .B(n6763), .Y(n1153) );
  OAI21X1 U2176 ( .A(n6486), .B(n6761), .C(n1154), .Y(n3565) );
  NAND2X1 U2177 ( .A(\Mem[39][31] ), .B(n6763), .Y(n1154) );
  NAND2X1 U2178 ( .A(n7011), .B(n7021), .Y(n1122) );
  NAND3X1 U2180 ( .A(n7015), .B(n7014), .C(n80), .Y(n1155) );
  OAI21X1 U2181 ( .A(n6606), .B(n6755), .C(n1158), .Y(n3566) );
  NAND2X1 U2182 ( .A(\Mem[40][0] ), .B(n6758), .Y(n1158) );
  OAI21X1 U2183 ( .A(n6551), .B(n6754), .C(n1159), .Y(n3567) );
  NAND2X1 U2184 ( .A(\Mem[40][1] ), .B(n6758), .Y(n1159) );
  OAI21X1 U2185 ( .A(n6496), .B(n6754), .C(n1160), .Y(n3568) );
  NAND2X1 U2186 ( .A(\Mem[40][2] ), .B(n6758), .Y(n1160) );
  OAI21X1 U2187 ( .A(n6481), .B(n6754), .C(n1161), .Y(n3569) );
  NAND2X1 U2188 ( .A(\Mem[40][3] ), .B(n6757), .Y(n1161) );
  OAI21X1 U2189 ( .A(n6476), .B(n6754), .C(n1162), .Y(n3570) );
  NAND2X1 U2190 ( .A(\Mem[40][4] ), .B(n6758), .Y(n1162) );
  OAI21X1 U2191 ( .A(n6471), .B(n6754), .C(n1163), .Y(n3571) );
  NAND2X1 U2192 ( .A(\Mem[40][5] ), .B(n6757), .Y(n1163) );
  OAI21X1 U2193 ( .A(n6466), .B(n6754), .C(n1164), .Y(n3572) );
  NAND2X1 U2194 ( .A(\Mem[40][6] ), .B(n6757), .Y(n1164) );
  OAI21X1 U2195 ( .A(n6461), .B(n6754), .C(n1165), .Y(n3573) );
  NAND2X1 U2196 ( .A(\Mem[40][7] ), .B(n6757), .Y(n1165) );
  OAI21X1 U2197 ( .A(n6456), .B(n6754), .C(n1166), .Y(n3574) );
  NAND2X1 U2198 ( .A(\Mem[40][8] ), .B(n6757), .Y(n1166) );
  OAI21X1 U2199 ( .A(n6451), .B(n6754), .C(n1167), .Y(n3575) );
  NAND2X1 U2200 ( .A(\Mem[40][9] ), .B(n6757), .Y(n1167) );
  OAI21X1 U2201 ( .A(n6601), .B(n6754), .C(n1168), .Y(n3576) );
  NAND2X1 U2202 ( .A(\Mem[40][10] ), .B(n6757), .Y(n1168) );
  OAI21X1 U2203 ( .A(n6596), .B(n6754), .C(n1169), .Y(n3577) );
  NAND2X1 U2204 ( .A(\Mem[40][11] ), .B(n6757), .Y(n1169) );
  OAI21X1 U2205 ( .A(n6591), .B(n6754), .C(n1170), .Y(n3578) );
  NAND2X1 U2206 ( .A(\Mem[40][12] ), .B(n6757), .Y(n1170) );
  OAI21X1 U2207 ( .A(n6586), .B(n6755), .C(n1171), .Y(n3579) );
  NAND2X1 U2208 ( .A(\Mem[40][13] ), .B(n6757), .Y(n1171) );
  OAI21X1 U2209 ( .A(n6581), .B(n6755), .C(n1172), .Y(n3580) );
  NAND2X1 U2210 ( .A(\Mem[40][14] ), .B(n6757), .Y(n1172) );
  OAI21X1 U2211 ( .A(n6576), .B(n6755), .C(n1173), .Y(n3581) );
  NAND2X1 U2212 ( .A(\Mem[40][15] ), .B(n6756), .Y(n1173) );
  OAI21X1 U2213 ( .A(n6571), .B(n6755), .C(n1174), .Y(n3582) );
  NAND2X1 U2214 ( .A(\Mem[40][16] ), .B(n6757), .Y(n1174) );
  OAI21X1 U2215 ( .A(n6566), .B(n6755), .C(n1175), .Y(n3583) );
  NAND2X1 U2216 ( .A(\Mem[40][17] ), .B(n6756), .Y(n1175) );
  OAI21X1 U2217 ( .A(n6561), .B(n6755), .C(n1176), .Y(n3584) );
  NAND2X1 U2218 ( .A(\Mem[40][18] ), .B(n6756), .Y(n1176) );
  OAI21X1 U2219 ( .A(n6556), .B(n6755), .C(n1177), .Y(n3585) );
  NAND2X1 U2220 ( .A(\Mem[40][19] ), .B(n6756), .Y(n1177) );
  OAI21X1 U2221 ( .A(n6546), .B(n6755), .C(n1178), .Y(n3586) );
  NAND2X1 U2222 ( .A(\Mem[40][20] ), .B(n6756), .Y(n1178) );
  OAI21X1 U2223 ( .A(n6541), .B(n6755), .C(n1179), .Y(n3587) );
  NAND2X1 U2224 ( .A(\Mem[40][21] ), .B(n6756), .Y(n1179) );
  OAI21X1 U2225 ( .A(n6536), .B(n6755), .C(n1180), .Y(n3588) );
  NAND2X1 U2226 ( .A(\Mem[40][22] ), .B(n6757), .Y(n1180) );
  OAI21X1 U2227 ( .A(n6531), .B(n6756), .C(n1181), .Y(n3589) );
  NAND2X1 U2228 ( .A(\Mem[40][23] ), .B(n6756), .Y(n1181) );
  OAI21X1 U2229 ( .A(n6526), .B(n6755), .C(n1182), .Y(n3590) );
  NAND2X1 U2230 ( .A(\Mem[40][24] ), .B(n6757), .Y(n1182) );
  OAI21X1 U2231 ( .A(n6521), .B(n6756), .C(n1183), .Y(n3591) );
  NAND2X1 U2232 ( .A(\Mem[40][25] ), .B(n6757), .Y(n1183) );
  OAI21X1 U2233 ( .A(n6516), .B(n6756), .C(n1184), .Y(n3592) );
  NAND2X1 U2234 ( .A(\Mem[40][26] ), .B(n6757), .Y(n1184) );
  OAI21X1 U2235 ( .A(n6511), .B(n6756), .C(n1185), .Y(n3593) );
  NAND2X1 U2236 ( .A(\Mem[40][27] ), .B(n6757), .Y(n1185) );
  OAI21X1 U2237 ( .A(n6506), .B(n6756), .C(n1186), .Y(n3594) );
  NAND2X1 U2238 ( .A(\Mem[40][28] ), .B(n6757), .Y(n1186) );
  OAI21X1 U2239 ( .A(n6501), .B(n6756), .C(n1187), .Y(n3595) );
  NAND2X1 U2240 ( .A(\Mem[40][29] ), .B(n6757), .Y(n1187) );
  OAI21X1 U2241 ( .A(n6491), .B(n6756), .C(n1188), .Y(n3596) );
  NAND2X1 U2242 ( .A(\Mem[40][30] ), .B(n6758), .Y(n1188) );
  OAI21X1 U2243 ( .A(n6486), .B(n6756), .C(n1189), .Y(n3597) );
  NAND2X1 U2244 ( .A(\Mem[40][31] ), .B(n6758), .Y(n1189) );
  NAND2X1 U2245 ( .A(n7010), .B(n7016), .Y(n1157) );
  OAI21X1 U2246 ( .A(n6606), .B(n6750), .C(n1192), .Y(n3598) );
  NAND2X1 U2247 ( .A(\Mem[41][0] ), .B(n6753), .Y(n1192) );
  OAI21X1 U2248 ( .A(n6551), .B(n6749), .C(n1193), .Y(n3599) );
  NAND2X1 U2249 ( .A(\Mem[41][1] ), .B(n6753), .Y(n1193) );
  OAI21X1 U2250 ( .A(n6496), .B(n6749), .C(n1194), .Y(n3600) );
  NAND2X1 U2251 ( .A(\Mem[41][2] ), .B(n6753), .Y(n1194) );
  OAI21X1 U2252 ( .A(n6481), .B(n6749), .C(n1195), .Y(n3601) );
  NAND2X1 U2253 ( .A(\Mem[41][3] ), .B(n6752), .Y(n1195) );
  OAI21X1 U2254 ( .A(n6476), .B(n6749), .C(n1196), .Y(n3602) );
  NAND2X1 U2255 ( .A(\Mem[41][4] ), .B(n6753), .Y(n1196) );
  OAI21X1 U2256 ( .A(n6471), .B(n6749), .C(n1197), .Y(n3603) );
  NAND2X1 U2257 ( .A(\Mem[41][5] ), .B(n6752), .Y(n1197) );
  OAI21X1 U2258 ( .A(n6466), .B(n6749), .C(n1198), .Y(n3604) );
  NAND2X1 U2259 ( .A(\Mem[41][6] ), .B(n6752), .Y(n1198) );
  OAI21X1 U2260 ( .A(n6461), .B(n6749), .C(n1199), .Y(n3605) );
  NAND2X1 U2261 ( .A(\Mem[41][7] ), .B(n6752), .Y(n1199) );
  OAI21X1 U2262 ( .A(n6456), .B(n6749), .C(n1200), .Y(n3606) );
  NAND2X1 U2263 ( .A(\Mem[41][8] ), .B(n6752), .Y(n1200) );
  OAI21X1 U2264 ( .A(n6451), .B(n6749), .C(n1201), .Y(n3607) );
  NAND2X1 U2265 ( .A(\Mem[41][9] ), .B(n6752), .Y(n1201) );
  OAI21X1 U2266 ( .A(n6601), .B(n6749), .C(n1202), .Y(n3608) );
  NAND2X1 U2267 ( .A(\Mem[41][10] ), .B(n6752), .Y(n1202) );
  OAI21X1 U2268 ( .A(n6596), .B(n6749), .C(n1203), .Y(n3609) );
  NAND2X1 U2269 ( .A(\Mem[41][11] ), .B(n6752), .Y(n1203) );
  OAI21X1 U2270 ( .A(n6591), .B(n6749), .C(n1204), .Y(n3610) );
  NAND2X1 U2271 ( .A(\Mem[41][12] ), .B(n6752), .Y(n1204) );
  OAI21X1 U2272 ( .A(n6586), .B(n6750), .C(n1205), .Y(n3611) );
  NAND2X1 U2273 ( .A(\Mem[41][13] ), .B(n6752), .Y(n1205) );
  OAI21X1 U2274 ( .A(n6581), .B(n6750), .C(n1206), .Y(n3612) );
  NAND2X1 U2275 ( .A(\Mem[41][14] ), .B(n6752), .Y(n1206) );
  OAI21X1 U2276 ( .A(n6576), .B(n6750), .C(n1207), .Y(n3613) );
  NAND2X1 U2277 ( .A(\Mem[41][15] ), .B(n6751), .Y(n1207) );
  OAI21X1 U2278 ( .A(n6571), .B(n6750), .C(n1208), .Y(n3614) );
  NAND2X1 U2279 ( .A(\Mem[41][16] ), .B(n6752), .Y(n1208) );
  OAI21X1 U2280 ( .A(n6566), .B(n6750), .C(n1209), .Y(n3615) );
  NAND2X1 U2281 ( .A(\Mem[41][17] ), .B(n6751), .Y(n1209) );
  OAI21X1 U2282 ( .A(n6561), .B(n6750), .C(n1210), .Y(n3616) );
  NAND2X1 U2283 ( .A(\Mem[41][18] ), .B(n6751), .Y(n1210) );
  OAI21X1 U2284 ( .A(n6556), .B(n6750), .C(n1211), .Y(n3617) );
  NAND2X1 U2285 ( .A(\Mem[41][19] ), .B(n6751), .Y(n1211) );
  OAI21X1 U2286 ( .A(n6546), .B(n6750), .C(n1212), .Y(n3618) );
  NAND2X1 U2287 ( .A(\Mem[41][20] ), .B(n6751), .Y(n1212) );
  OAI21X1 U2288 ( .A(n6541), .B(n6750), .C(n1213), .Y(n3619) );
  NAND2X1 U2289 ( .A(\Mem[41][21] ), .B(n6751), .Y(n1213) );
  OAI21X1 U2290 ( .A(n6536), .B(n6750), .C(n1214), .Y(n3620) );
  NAND2X1 U2291 ( .A(\Mem[41][22] ), .B(n6752), .Y(n1214) );
  OAI21X1 U2292 ( .A(n6531), .B(n6751), .C(n1215), .Y(n3621) );
  NAND2X1 U2293 ( .A(\Mem[41][23] ), .B(n6751), .Y(n1215) );
  OAI21X1 U2294 ( .A(n6526), .B(n6750), .C(n1216), .Y(n3622) );
  NAND2X1 U2295 ( .A(\Mem[41][24] ), .B(n6752), .Y(n1216) );
  OAI21X1 U2296 ( .A(n6521), .B(n6751), .C(n1217), .Y(n3623) );
  NAND2X1 U2297 ( .A(\Mem[41][25] ), .B(n6752), .Y(n1217) );
  OAI21X1 U2298 ( .A(n6516), .B(n6751), .C(n1218), .Y(n3624) );
  NAND2X1 U2299 ( .A(\Mem[41][26] ), .B(n6752), .Y(n1218) );
  OAI21X1 U2300 ( .A(n6511), .B(n6751), .C(n1219), .Y(n3625) );
  NAND2X1 U2301 ( .A(\Mem[41][27] ), .B(n6752), .Y(n1219) );
  OAI21X1 U2302 ( .A(n6506), .B(n6751), .C(n1220), .Y(n3626) );
  NAND2X1 U2303 ( .A(\Mem[41][28] ), .B(n6752), .Y(n1220) );
  OAI21X1 U2304 ( .A(n6501), .B(n6751), .C(n1221), .Y(n3627) );
  NAND2X1 U2305 ( .A(\Mem[41][29] ), .B(n6752), .Y(n1221) );
  OAI21X1 U2306 ( .A(n6491), .B(n6751), .C(n1222), .Y(n3628) );
  NAND2X1 U2307 ( .A(\Mem[41][30] ), .B(n6753), .Y(n1222) );
  OAI21X1 U2308 ( .A(n6486), .B(n6751), .C(n1223), .Y(n3629) );
  NAND2X1 U2309 ( .A(\Mem[41][31] ), .B(n6753), .Y(n1223) );
  NAND2X1 U2310 ( .A(n7010), .B(n7017), .Y(n1191) );
  OAI21X1 U2311 ( .A(n6606), .B(n6745), .C(n1225), .Y(n3630) );
  NAND2X1 U2312 ( .A(\Mem[42][0] ), .B(n6748), .Y(n1225) );
  OAI21X1 U2313 ( .A(n6551), .B(n6744), .C(n1226), .Y(n3631) );
  NAND2X1 U2314 ( .A(\Mem[42][1] ), .B(n6748), .Y(n1226) );
  OAI21X1 U2315 ( .A(n6496), .B(n6744), .C(n1227), .Y(n3632) );
  NAND2X1 U2316 ( .A(\Mem[42][2] ), .B(n6748), .Y(n1227) );
  OAI21X1 U2317 ( .A(n6481), .B(n6744), .C(n1228), .Y(n3633) );
  NAND2X1 U2318 ( .A(\Mem[42][3] ), .B(n6747), .Y(n1228) );
  OAI21X1 U2319 ( .A(n6476), .B(n6744), .C(n1229), .Y(n3634) );
  NAND2X1 U2320 ( .A(\Mem[42][4] ), .B(n6748), .Y(n1229) );
  OAI21X1 U2321 ( .A(n6471), .B(n6744), .C(n1230), .Y(n3635) );
  NAND2X1 U2322 ( .A(\Mem[42][5] ), .B(n6747), .Y(n1230) );
  OAI21X1 U2323 ( .A(n6466), .B(n6744), .C(n1231), .Y(n3636) );
  NAND2X1 U2324 ( .A(\Mem[42][6] ), .B(n6747), .Y(n1231) );
  OAI21X1 U2325 ( .A(n6461), .B(n6744), .C(n1232), .Y(n3637) );
  NAND2X1 U2326 ( .A(\Mem[42][7] ), .B(n6747), .Y(n1232) );
  OAI21X1 U2327 ( .A(n6456), .B(n6744), .C(n1233), .Y(n3638) );
  NAND2X1 U2328 ( .A(\Mem[42][8] ), .B(n6747), .Y(n1233) );
  OAI21X1 U2329 ( .A(n6451), .B(n6744), .C(n1234), .Y(n3639) );
  NAND2X1 U2330 ( .A(\Mem[42][9] ), .B(n6747), .Y(n1234) );
  OAI21X1 U2331 ( .A(n6601), .B(n6744), .C(n1235), .Y(n3640) );
  NAND2X1 U2332 ( .A(\Mem[42][10] ), .B(n6747), .Y(n1235) );
  OAI21X1 U2333 ( .A(n6596), .B(n6744), .C(n1236), .Y(n3641) );
  NAND2X1 U2334 ( .A(\Mem[42][11] ), .B(n6747), .Y(n1236) );
  OAI21X1 U2335 ( .A(n6591), .B(n6744), .C(n1237), .Y(n3642) );
  NAND2X1 U2336 ( .A(\Mem[42][12] ), .B(n6747), .Y(n1237) );
  OAI21X1 U2337 ( .A(n6586), .B(n6745), .C(n1238), .Y(n3643) );
  NAND2X1 U2338 ( .A(\Mem[42][13] ), .B(n6747), .Y(n1238) );
  OAI21X1 U2339 ( .A(n6581), .B(n6745), .C(n1239), .Y(n3644) );
  NAND2X1 U2340 ( .A(\Mem[42][14] ), .B(n6747), .Y(n1239) );
  OAI21X1 U2341 ( .A(n6576), .B(n6745), .C(n1240), .Y(n3645) );
  NAND2X1 U2342 ( .A(\Mem[42][15] ), .B(n6746), .Y(n1240) );
  OAI21X1 U2343 ( .A(n6571), .B(n6745), .C(n1241), .Y(n3646) );
  NAND2X1 U2344 ( .A(\Mem[42][16] ), .B(n6747), .Y(n1241) );
  OAI21X1 U2345 ( .A(n6566), .B(n6745), .C(n1242), .Y(n3647) );
  NAND2X1 U2346 ( .A(\Mem[42][17] ), .B(n6746), .Y(n1242) );
  OAI21X1 U2347 ( .A(n6561), .B(n6745), .C(n1243), .Y(n3648) );
  NAND2X1 U2348 ( .A(\Mem[42][18] ), .B(n6746), .Y(n1243) );
  OAI21X1 U2349 ( .A(n6556), .B(n6745), .C(n1244), .Y(n3649) );
  NAND2X1 U2350 ( .A(\Mem[42][19] ), .B(n6746), .Y(n1244) );
  OAI21X1 U2351 ( .A(n6546), .B(n6745), .C(n1245), .Y(n3650) );
  NAND2X1 U2352 ( .A(\Mem[42][20] ), .B(n6746), .Y(n1245) );
  OAI21X1 U2353 ( .A(n6541), .B(n6745), .C(n1246), .Y(n3651) );
  NAND2X1 U2354 ( .A(\Mem[42][21] ), .B(n6746), .Y(n1246) );
  OAI21X1 U2355 ( .A(n6536), .B(n6745), .C(n1247), .Y(n3652) );
  NAND2X1 U2356 ( .A(\Mem[42][22] ), .B(n6747), .Y(n1247) );
  OAI21X1 U2357 ( .A(n6531), .B(n6746), .C(n1248), .Y(n3653) );
  NAND2X1 U2358 ( .A(\Mem[42][23] ), .B(n6746), .Y(n1248) );
  OAI21X1 U2359 ( .A(n6526), .B(n6745), .C(n1249), .Y(n3654) );
  NAND2X1 U2360 ( .A(\Mem[42][24] ), .B(n6747), .Y(n1249) );
  OAI21X1 U2361 ( .A(n6521), .B(n6746), .C(n1250), .Y(n3655) );
  NAND2X1 U2362 ( .A(\Mem[42][25] ), .B(n6747), .Y(n1250) );
  OAI21X1 U2363 ( .A(n6516), .B(n6746), .C(n1251), .Y(n3656) );
  NAND2X1 U2364 ( .A(\Mem[42][26] ), .B(n6747), .Y(n1251) );
  OAI21X1 U2365 ( .A(n6511), .B(n6746), .C(n1252), .Y(n3657) );
  NAND2X1 U2366 ( .A(\Mem[42][27] ), .B(n6747), .Y(n1252) );
  OAI21X1 U2367 ( .A(n6506), .B(n6746), .C(n1253), .Y(n3658) );
  NAND2X1 U2368 ( .A(\Mem[42][28] ), .B(n6747), .Y(n1253) );
  OAI21X1 U2369 ( .A(n6501), .B(n6746), .C(n1254), .Y(n3659) );
  NAND2X1 U2370 ( .A(\Mem[42][29] ), .B(n6747), .Y(n1254) );
  OAI21X1 U2371 ( .A(n6491), .B(n6746), .C(n1255), .Y(n3660) );
  NAND2X1 U2372 ( .A(\Mem[42][30] ), .B(n6748), .Y(n1255) );
  OAI21X1 U2373 ( .A(n6486), .B(n6746), .C(n1256), .Y(n3661) );
  NAND2X1 U2374 ( .A(\Mem[42][31] ), .B(n6748), .Y(n1256) );
  NAND2X1 U2375 ( .A(n7010), .B(n7018), .Y(n1224) );
  OAI21X1 U2376 ( .A(n6606), .B(n6740), .C(n1258), .Y(n3662) );
  NAND2X1 U2377 ( .A(\Mem[43][0] ), .B(n6743), .Y(n1258) );
  OAI21X1 U2378 ( .A(n6551), .B(n6739), .C(n1259), .Y(n3663) );
  NAND2X1 U2379 ( .A(\Mem[43][1] ), .B(n6743), .Y(n1259) );
  OAI21X1 U2380 ( .A(n6496), .B(n6739), .C(n1260), .Y(n3664) );
  NAND2X1 U2381 ( .A(\Mem[43][2] ), .B(n6743), .Y(n1260) );
  OAI21X1 U2382 ( .A(n6481), .B(n6739), .C(n1261), .Y(n3665) );
  NAND2X1 U2383 ( .A(\Mem[43][3] ), .B(n6742), .Y(n1261) );
  OAI21X1 U2384 ( .A(n6476), .B(n6739), .C(n1262), .Y(n3666) );
  NAND2X1 U2385 ( .A(\Mem[43][4] ), .B(n6743), .Y(n1262) );
  OAI21X1 U2386 ( .A(n6471), .B(n6739), .C(n1263), .Y(n3667) );
  NAND2X1 U2387 ( .A(\Mem[43][5] ), .B(n6742), .Y(n1263) );
  OAI21X1 U2388 ( .A(n6466), .B(n6739), .C(n1264), .Y(n3668) );
  NAND2X1 U2389 ( .A(\Mem[43][6] ), .B(n6742), .Y(n1264) );
  OAI21X1 U2390 ( .A(n6461), .B(n6739), .C(n1265), .Y(n3669) );
  NAND2X1 U2391 ( .A(\Mem[43][7] ), .B(n6742), .Y(n1265) );
  OAI21X1 U2392 ( .A(n6456), .B(n6739), .C(n1266), .Y(n3670) );
  NAND2X1 U2393 ( .A(\Mem[43][8] ), .B(n6742), .Y(n1266) );
  OAI21X1 U2394 ( .A(n6451), .B(n6739), .C(n1267), .Y(n3671) );
  NAND2X1 U2395 ( .A(\Mem[43][9] ), .B(n6742), .Y(n1267) );
  OAI21X1 U2396 ( .A(n6601), .B(n6739), .C(n1268), .Y(n3672) );
  NAND2X1 U2397 ( .A(\Mem[43][10] ), .B(n6742), .Y(n1268) );
  OAI21X1 U2398 ( .A(n6596), .B(n6739), .C(n1269), .Y(n3673) );
  NAND2X1 U2399 ( .A(\Mem[43][11] ), .B(n6742), .Y(n1269) );
  OAI21X1 U2400 ( .A(n6591), .B(n6739), .C(n1270), .Y(n3674) );
  NAND2X1 U2401 ( .A(\Mem[43][12] ), .B(n6742), .Y(n1270) );
  OAI21X1 U2402 ( .A(n6586), .B(n6740), .C(n1271), .Y(n3675) );
  NAND2X1 U2403 ( .A(\Mem[43][13] ), .B(n6742), .Y(n1271) );
  OAI21X1 U2404 ( .A(n6581), .B(n6740), .C(n1272), .Y(n3676) );
  NAND2X1 U2405 ( .A(\Mem[43][14] ), .B(n6742), .Y(n1272) );
  OAI21X1 U2406 ( .A(n6576), .B(n6740), .C(n1273), .Y(n3677) );
  NAND2X1 U2407 ( .A(\Mem[43][15] ), .B(n6741), .Y(n1273) );
  OAI21X1 U2408 ( .A(n6571), .B(n6740), .C(n1274), .Y(n3678) );
  NAND2X1 U2409 ( .A(\Mem[43][16] ), .B(n6742), .Y(n1274) );
  OAI21X1 U2410 ( .A(n6566), .B(n6740), .C(n1275), .Y(n3679) );
  NAND2X1 U2411 ( .A(\Mem[43][17] ), .B(n6741), .Y(n1275) );
  OAI21X1 U2412 ( .A(n6561), .B(n6740), .C(n1276), .Y(n3680) );
  NAND2X1 U2413 ( .A(\Mem[43][18] ), .B(n6741), .Y(n1276) );
  OAI21X1 U2414 ( .A(n6556), .B(n6740), .C(n1277), .Y(n3681) );
  NAND2X1 U2415 ( .A(\Mem[43][19] ), .B(n6741), .Y(n1277) );
  OAI21X1 U2416 ( .A(n6546), .B(n6740), .C(n1278), .Y(n3682) );
  NAND2X1 U2417 ( .A(\Mem[43][20] ), .B(n6741), .Y(n1278) );
  OAI21X1 U2418 ( .A(n6541), .B(n6740), .C(n1279), .Y(n3683) );
  NAND2X1 U2419 ( .A(\Mem[43][21] ), .B(n6741), .Y(n1279) );
  OAI21X1 U2420 ( .A(n6536), .B(n6740), .C(n1280), .Y(n3684) );
  NAND2X1 U2421 ( .A(\Mem[43][22] ), .B(n6742), .Y(n1280) );
  OAI21X1 U2422 ( .A(n6531), .B(n6741), .C(n1281), .Y(n3685) );
  NAND2X1 U2423 ( .A(\Mem[43][23] ), .B(n6741), .Y(n1281) );
  OAI21X1 U2424 ( .A(n6526), .B(n6740), .C(n1282), .Y(n3686) );
  NAND2X1 U2425 ( .A(\Mem[43][24] ), .B(n6742), .Y(n1282) );
  OAI21X1 U2426 ( .A(n6521), .B(n6741), .C(n1283), .Y(n3687) );
  NAND2X1 U2427 ( .A(\Mem[43][25] ), .B(n6742), .Y(n1283) );
  OAI21X1 U2428 ( .A(n6516), .B(n6741), .C(n1284), .Y(n3688) );
  NAND2X1 U2429 ( .A(\Mem[43][26] ), .B(n6742), .Y(n1284) );
  OAI21X1 U2430 ( .A(n6511), .B(n6741), .C(n1285), .Y(n3689) );
  NAND2X1 U2431 ( .A(\Mem[43][27] ), .B(n6742), .Y(n1285) );
  OAI21X1 U2432 ( .A(n6506), .B(n6741), .C(n1286), .Y(n3690) );
  NAND2X1 U2433 ( .A(\Mem[43][28] ), .B(n6742), .Y(n1286) );
  OAI21X1 U2434 ( .A(n6501), .B(n6741), .C(n1287), .Y(n3691) );
  NAND2X1 U2435 ( .A(\Mem[43][29] ), .B(n6742), .Y(n1287) );
  OAI21X1 U2436 ( .A(n6491), .B(n6741), .C(n1288), .Y(n3692) );
  NAND2X1 U2437 ( .A(\Mem[43][30] ), .B(n6743), .Y(n1288) );
  OAI21X1 U2438 ( .A(n6486), .B(n6741), .C(n1289), .Y(n3693) );
  NAND2X1 U2439 ( .A(\Mem[43][31] ), .B(n6743), .Y(n1289) );
  NAND2X1 U2440 ( .A(n7010), .B(n7019), .Y(n1257) );
  OAI21X1 U2441 ( .A(n6607), .B(n6735), .C(n1291), .Y(n3694) );
  NAND2X1 U2442 ( .A(\Mem[44][0] ), .B(n6738), .Y(n1291) );
  OAI21X1 U2443 ( .A(n6552), .B(n6734), .C(n1292), .Y(n3695) );
  NAND2X1 U2444 ( .A(\Mem[44][1] ), .B(n6738), .Y(n1292) );
  OAI21X1 U2445 ( .A(n6497), .B(n6734), .C(n1293), .Y(n3696) );
  NAND2X1 U2446 ( .A(\Mem[44][2] ), .B(n6738), .Y(n1293) );
  OAI21X1 U2447 ( .A(n6482), .B(n6734), .C(n1294), .Y(n3697) );
  NAND2X1 U2448 ( .A(\Mem[44][3] ), .B(n6737), .Y(n1294) );
  OAI21X1 U2449 ( .A(n6477), .B(n6734), .C(n1295), .Y(n3698) );
  NAND2X1 U2450 ( .A(\Mem[44][4] ), .B(n6738), .Y(n1295) );
  OAI21X1 U2451 ( .A(n6472), .B(n6734), .C(n1296), .Y(n3699) );
  NAND2X1 U2452 ( .A(\Mem[44][5] ), .B(n6737), .Y(n1296) );
  OAI21X1 U2453 ( .A(n6467), .B(n6734), .C(n1297), .Y(n3700) );
  NAND2X1 U2454 ( .A(\Mem[44][6] ), .B(n6737), .Y(n1297) );
  OAI21X1 U2455 ( .A(n6462), .B(n6734), .C(n1298), .Y(n3701) );
  NAND2X1 U2456 ( .A(\Mem[44][7] ), .B(n6737), .Y(n1298) );
  OAI21X1 U2457 ( .A(n6457), .B(n6734), .C(n1299), .Y(n3702) );
  NAND2X1 U2458 ( .A(\Mem[44][8] ), .B(n6737), .Y(n1299) );
  OAI21X1 U2459 ( .A(n6452), .B(n6734), .C(n1300), .Y(n3703) );
  NAND2X1 U2460 ( .A(\Mem[44][9] ), .B(n6737), .Y(n1300) );
  OAI21X1 U2461 ( .A(n6602), .B(n6734), .C(n1301), .Y(n3704) );
  NAND2X1 U2462 ( .A(\Mem[44][10] ), .B(n6737), .Y(n1301) );
  OAI21X1 U2463 ( .A(n6597), .B(n6734), .C(n1302), .Y(n3705) );
  NAND2X1 U2464 ( .A(\Mem[44][11] ), .B(n6737), .Y(n1302) );
  OAI21X1 U2465 ( .A(n6592), .B(n6734), .C(n1303), .Y(n3706) );
  NAND2X1 U2466 ( .A(\Mem[44][12] ), .B(n6737), .Y(n1303) );
  OAI21X1 U2467 ( .A(n6587), .B(n6735), .C(n1304), .Y(n3707) );
  NAND2X1 U2468 ( .A(\Mem[44][13] ), .B(n6737), .Y(n1304) );
  OAI21X1 U2469 ( .A(n6582), .B(n6735), .C(n1305), .Y(n3708) );
  NAND2X1 U2470 ( .A(\Mem[44][14] ), .B(n6737), .Y(n1305) );
  OAI21X1 U2471 ( .A(n6577), .B(n6735), .C(n1306), .Y(n3709) );
  NAND2X1 U2472 ( .A(\Mem[44][15] ), .B(n6736), .Y(n1306) );
  OAI21X1 U2473 ( .A(n6572), .B(n6735), .C(n1307), .Y(n3710) );
  NAND2X1 U2474 ( .A(\Mem[44][16] ), .B(n6737), .Y(n1307) );
  OAI21X1 U2475 ( .A(n6567), .B(n6735), .C(n1308), .Y(n3711) );
  NAND2X1 U2476 ( .A(\Mem[44][17] ), .B(n6736), .Y(n1308) );
  OAI21X1 U2477 ( .A(n6562), .B(n6735), .C(n1309), .Y(n3712) );
  NAND2X1 U2478 ( .A(\Mem[44][18] ), .B(n6736), .Y(n1309) );
  OAI21X1 U2479 ( .A(n6556), .B(n6735), .C(n1310), .Y(n3713) );
  NAND2X1 U2480 ( .A(\Mem[44][19] ), .B(n6736), .Y(n1310) );
  OAI21X1 U2481 ( .A(n6546), .B(n6735), .C(n1311), .Y(n3714) );
  NAND2X1 U2482 ( .A(\Mem[44][20] ), .B(n6736), .Y(n1311) );
  OAI21X1 U2483 ( .A(n6541), .B(n6735), .C(n1312), .Y(n3715) );
  NAND2X1 U2484 ( .A(\Mem[44][21] ), .B(n6736), .Y(n1312) );
  OAI21X1 U2485 ( .A(n6536), .B(n6735), .C(n1313), .Y(n3716) );
  NAND2X1 U2486 ( .A(\Mem[44][22] ), .B(n6737), .Y(n1313) );
  OAI21X1 U2487 ( .A(n6531), .B(n6736), .C(n1314), .Y(n3717) );
  NAND2X1 U2488 ( .A(\Mem[44][23] ), .B(n6736), .Y(n1314) );
  OAI21X1 U2489 ( .A(n6526), .B(n6735), .C(n1315), .Y(n3718) );
  NAND2X1 U2490 ( .A(\Mem[44][24] ), .B(n6737), .Y(n1315) );
  OAI21X1 U2491 ( .A(n6521), .B(n6736), .C(n1316), .Y(n3719) );
  NAND2X1 U2492 ( .A(\Mem[44][25] ), .B(n6737), .Y(n1316) );
  OAI21X1 U2493 ( .A(n6516), .B(n6736), .C(n1317), .Y(n3720) );
  NAND2X1 U2494 ( .A(\Mem[44][26] ), .B(n6737), .Y(n1317) );
  OAI21X1 U2495 ( .A(n6511), .B(n6736), .C(n1318), .Y(n3721) );
  NAND2X1 U2496 ( .A(\Mem[44][27] ), .B(n6737), .Y(n1318) );
  OAI21X1 U2497 ( .A(n6506), .B(n6736), .C(n1319), .Y(n3722) );
  NAND2X1 U2498 ( .A(\Mem[44][28] ), .B(n6737), .Y(n1319) );
  OAI21X1 U2499 ( .A(n6501), .B(n6736), .C(n1320), .Y(n3723) );
  NAND2X1 U2500 ( .A(\Mem[44][29] ), .B(n6737), .Y(n1320) );
  OAI21X1 U2501 ( .A(n6491), .B(n6736), .C(n1321), .Y(n3724) );
  NAND2X1 U2502 ( .A(\Mem[44][30] ), .B(n6738), .Y(n1321) );
  OAI21X1 U2503 ( .A(n6486), .B(n6736), .C(n1322), .Y(n3725) );
  NAND2X1 U2504 ( .A(\Mem[44][31] ), .B(n6738), .Y(n1322) );
  NAND2X1 U2505 ( .A(n7010), .B(n7022), .Y(n1290) );
  OAI21X1 U2506 ( .A(n6607), .B(n6730), .C(n1324), .Y(n3726) );
  NAND2X1 U2507 ( .A(\Mem[45][0] ), .B(n6733), .Y(n1324) );
  OAI21X1 U2508 ( .A(n6552), .B(n6729), .C(n1325), .Y(n3727) );
  NAND2X1 U2509 ( .A(\Mem[45][1] ), .B(n6733), .Y(n1325) );
  OAI21X1 U2510 ( .A(n6497), .B(n6729), .C(n1326), .Y(n3728) );
  NAND2X1 U2511 ( .A(\Mem[45][2] ), .B(n6733), .Y(n1326) );
  OAI21X1 U2512 ( .A(n6482), .B(n6729), .C(n1327), .Y(n3729) );
  NAND2X1 U2513 ( .A(\Mem[45][3] ), .B(n6732), .Y(n1327) );
  OAI21X1 U2514 ( .A(n6477), .B(n6729), .C(n1328), .Y(n3730) );
  NAND2X1 U2515 ( .A(\Mem[45][4] ), .B(n6733), .Y(n1328) );
  OAI21X1 U2516 ( .A(n6472), .B(n6729), .C(n1329), .Y(n3731) );
  NAND2X1 U2517 ( .A(\Mem[45][5] ), .B(n6732), .Y(n1329) );
  OAI21X1 U2518 ( .A(n6467), .B(n6729), .C(n1330), .Y(n3732) );
  NAND2X1 U2519 ( .A(\Mem[45][6] ), .B(n6732), .Y(n1330) );
  OAI21X1 U2520 ( .A(n6462), .B(n6729), .C(n1331), .Y(n3733) );
  NAND2X1 U2521 ( .A(\Mem[45][7] ), .B(n6732), .Y(n1331) );
  OAI21X1 U2522 ( .A(n6457), .B(n6729), .C(n1332), .Y(n3734) );
  NAND2X1 U2523 ( .A(\Mem[45][8] ), .B(n6732), .Y(n1332) );
  OAI21X1 U2524 ( .A(n6452), .B(n6729), .C(n1333), .Y(n3735) );
  NAND2X1 U2525 ( .A(\Mem[45][9] ), .B(n6732), .Y(n1333) );
  OAI21X1 U2526 ( .A(n6602), .B(n6729), .C(n1334), .Y(n3736) );
  NAND2X1 U2527 ( .A(\Mem[45][10] ), .B(n6732), .Y(n1334) );
  OAI21X1 U2528 ( .A(n6597), .B(n6729), .C(n1335), .Y(n3737) );
  NAND2X1 U2529 ( .A(\Mem[45][11] ), .B(n6732), .Y(n1335) );
  OAI21X1 U2530 ( .A(n6592), .B(n6729), .C(n1336), .Y(n3738) );
  NAND2X1 U2531 ( .A(\Mem[45][12] ), .B(n6732), .Y(n1336) );
  OAI21X1 U2532 ( .A(n6587), .B(n6730), .C(n1337), .Y(n3739) );
  NAND2X1 U2533 ( .A(\Mem[45][13] ), .B(n6732), .Y(n1337) );
  OAI21X1 U2534 ( .A(n6582), .B(n6730), .C(n1338), .Y(n3740) );
  NAND2X1 U2535 ( .A(\Mem[45][14] ), .B(n6732), .Y(n1338) );
  OAI21X1 U2536 ( .A(n6577), .B(n6730), .C(n1339), .Y(n3741) );
  NAND2X1 U2537 ( .A(\Mem[45][15] ), .B(n6731), .Y(n1339) );
  OAI21X1 U2538 ( .A(n6572), .B(n6730), .C(n1340), .Y(n3742) );
  NAND2X1 U2539 ( .A(\Mem[45][16] ), .B(n6732), .Y(n1340) );
  OAI21X1 U2540 ( .A(n6567), .B(n6730), .C(n1341), .Y(n3743) );
  NAND2X1 U2541 ( .A(\Mem[45][17] ), .B(n6731), .Y(n1341) );
  OAI21X1 U2542 ( .A(n6562), .B(n6730), .C(n1342), .Y(n3744) );
  NAND2X1 U2543 ( .A(\Mem[45][18] ), .B(n6731), .Y(n1342) );
  OAI21X1 U2544 ( .A(n6557), .B(n6730), .C(n1343), .Y(n3745) );
  NAND2X1 U2545 ( .A(\Mem[45][19] ), .B(n6731), .Y(n1343) );
  OAI21X1 U2546 ( .A(n6547), .B(n6730), .C(n1344), .Y(n3746) );
  NAND2X1 U2547 ( .A(\Mem[45][20] ), .B(n6731), .Y(n1344) );
  OAI21X1 U2548 ( .A(n6542), .B(n6730), .C(n1345), .Y(n3747) );
  NAND2X1 U2549 ( .A(\Mem[45][21] ), .B(n6731), .Y(n1345) );
  OAI21X1 U2550 ( .A(n6537), .B(n6730), .C(n1346), .Y(n3748) );
  NAND2X1 U2551 ( .A(\Mem[45][22] ), .B(n6732), .Y(n1346) );
  OAI21X1 U2552 ( .A(n6532), .B(n6731), .C(n1347), .Y(n3749) );
  NAND2X1 U2553 ( .A(\Mem[45][23] ), .B(n6731), .Y(n1347) );
  OAI21X1 U2554 ( .A(n6527), .B(n6730), .C(n1348), .Y(n3750) );
  NAND2X1 U2555 ( .A(\Mem[45][24] ), .B(n6732), .Y(n1348) );
  OAI21X1 U2556 ( .A(n6522), .B(n6731), .C(n1349), .Y(n3751) );
  NAND2X1 U2557 ( .A(\Mem[45][25] ), .B(n6732), .Y(n1349) );
  OAI21X1 U2558 ( .A(n6517), .B(n6731), .C(n1350), .Y(n3752) );
  NAND2X1 U2559 ( .A(\Mem[45][26] ), .B(n6732), .Y(n1350) );
  OAI21X1 U2560 ( .A(n6512), .B(n6731), .C(n1351), .Y(n3753) );
  NAND2X1 U2561 ( .A(\Mem[45][27] ), .B(n6732), .Y(n1351) );
  OAI21X1 U2562 ( .A(n6507), .B(n6731), .C(n1352), .Y(n3754) );
  NAND2X1 U2563 ( .A(\Mem[45][28] ), .B(n6732), .Y(n1352) );
  OAI21X1 U2564 ( .A(n6502), .B(n6731), .C(n1353), .Y(n3755) );
  NAND2X1 U2565 ( .A(\Mem[45][29] ), .B(n6732), .Y(n1353) );
  OAI21X1 U2566 ( .A(n6492), .B(n6731), .C(n1354), .Y(n3756) );
  NAND2X1 U2567 ( .A(\Mem[45][30] ), .B(n6733), .Y(n1354) );
  OAI21X1 U2568 ( .A(n6487), .B(n6731), .C(n1355), .Y(n3757) );
  NAND2X1 U2569 ( .A(\Mem[45][31] ), .B(n6733), .Y(n1355) );
  NAND2X1 U2570 ( .A(n7010), .B(n7023), .Y(n1323) );
  OAI21X1 U2571 ( .A(n6607), .B(n6725), .C(n1357), .Y(n3758) );
  NAND2X1 U2572 ( .A(\Mem[46][0] ), .B(n6728), .Y(n1357) );
  OAI21X1 U2573 ( .A(n6552), .B(n6724), .C(n1358), .Y(n3759) );
  NAND2X1 U2574 ( .A(\Mem[46][1] ), .B(n6728), .Y(n1358) );
  OAI21X1 U2575 ( .A(n6497), .B(n6724), .C(n1359), .Y(n3760) );
  NAND2X1 U2576 ( .A(\Mem[46][2] ), .B(n6728), .Y(n1359) );
  OAI21X1 U2577 ( .A(n6482), .B(n6724), .C(n1360), .Y(n3761) );
  NAND2X1 U2578 ( .A(\Mem[46][3] ), .B(n6727), .Y(n1360) );
  OAI21X1 U2579 ( .A(n6477), .B(n6724), .C(n1361), .Y(n3762) );
  NAND2X1 U2580 ( .A(\Mem[46][4] ), .B(n6728), .Y(n1361) );
  OAI21X1 U2581 ( .A(n6472), .B(n6724), .C(n1362), .Y(n3763) );
  NAND2X1 U2582 ( .A(\Mem[46][5] ), .B(n6727), .Y(n1362) );
  OAI21X1 U2583 ( .A(n6467), .B(n6724), .C(n1363), .Y(n3764) );
  NAND2X1 U2584 ( .A(\Mem[46][6] ), .B(n6727), .Y(n1363) );
  OAI21X1 U2585 ( .A(n6462), .B(n6724), .C(n1364), .Y(n3765) );
  NAND2X1 U2586 ( .A(\Mem[46][7] ), .B(n6727), .Y(n1364) );
  OAI21X1 U2587 ( .A(n6457), .B(n6724), .C(n1365), .Y(n3766) );
  NAND2X1 U2588 ( .A(\Mem[46][8] ), .B(n6727), .Y(n1365) );
  OAI21X1 U2589 ( .A(n6452), .B(n6724), .C(n1366), .Y(n3767) );
  NAND2X1 U2590 ( .A(\Mem[46][9] ), .B(n6727), .Y(n1366) );
  OAI21X1 U2591 ( .A(n6602), .B(n6724), .C(n1367), .Y(n3768) );
  NAND2X1 U2592 ( .A(\Mem[46][10] ), .B(n6727), .Y(n1367) );
  OAI21X1 U2593 ( .A(n6597), .B(n6724), .C(n1368), .Y(n3769) );
  NAND2X1 U2594 ( .A(\Mem[46][11] ), .B(n6727), .Y(n1368) );
  OAI21X1 U2595 ( .A(n6592), .B(n6724), .C(n1369), .Y(n3770) );
  NAND2X1 U2596 ( .A(\Mem[46][12] ), .B(n6727), .Y(n1369) );
  OAI21X1 U2597 ( .A(n6587), .B(n6725), .C(n1370), .Y(n3771) );
  NAND2X1 U2598 ( .A(\Mem[46][13] ), .B(n6727), .Y(n1370) );
  OAI21X1 U2599 ( .A(n6582), .B(n6725), .C(n1371), .Y(n3772) );
  NAND2X1 U2600 ( .A(\Mem[46][14] ), .B(n6727), .Y(n1371) );
  OAI21X1 U2601 ( .A(n6577), .B(n6725), .C(n1372), .Y(n3773) );
  NAND2X1 U2602 ( .A(\Mem[46][15] ), .B(n6726), .Y(n1372) );
  OAI21X1 U2603 ( .A(n6572), .B(n6725), .C(n1373), .Y(n3774) );
  NAND2X1 U2604 ( .A(\Mem[46][16] ), .B(n6727), .Y(n1373) );
  OAI21X1 U2605 ( .A(n6567), .B(n6725), .C(n1374), .Y(n3775) );
  NAND2X1 U2606 ( .A(\Mem[46][17] ), .B(n6726), .Y(n1374) );
  OAI21X1 U2607 ( .A(n6562), .B(n6725), .C(n1375), .Y(n3776) );
  NAND2X1 U2608 ( .A(\Mem[46][18] ), .B(n6726), .Y(n1375) );
  OAI21X1 U2609 ( .A(n6557), .B(n6725), .C(n1376), .Y(n3777) );
  NAND2X1 U2610 ( .A(\Mem[46][19] ), .B(n6726), .Y(n1376) );
  OAI21X1 U2611 ( .A(n6547), .B(n6725), .C(n1377), .Y(n3778) );
  NAND2X1 U2612 ( .A(\Mem[46][20] ), .B(n6726), .Y(n1377) );
  OAI21X1 U2613 ( .A(n6542), .B(n6725), .C(n1378), .Y(n3779) );
  NAND2X1 U2614 ( .A(\Mem[46][21] ), .B(n6726), .Y(n1378) );
  OAI21X1 U2615 ( .A(n6537), .B(n6725), .C(n1379), .Y(n3780) );
  NAND2X1 U2616 ( .A(\Mem[46][22] ), .B(n6727), .Y(n1379) );
  OAI21X1 U2617 ( .A(n6532), .B(n6726), .C(n1380), .Y(n3781) );
  NAND2X1 U2618 ( .A(\Mem[46][23] ), .B(n6726), .Y(n1380) );
  OAI21X1 U2619 ( .A(n6527), .B(n6725), .C(n1381), .Y(n3782) );
  NAND2X1 U2620 ( .A(\Mem[46][24] ), .B(n6727), .Y(n1381) );
  OAI21X1 U2621 ( .A(n6522), .B(n6726), .C(n1382), .Y(n3783) );
  NAND2X1 U2622 ( .A(\Mem[46][25] ), .B(n6727), .Y(n1382) );
  OAI21X1 U2623 ( .A(n6517), .B(n6726), .C(n1383), .Y(n3784) );
  NAND2X1 U2624 ( .A(\Mem[46][26] ), .B(n6727), .Y(n1383) );
  OAI21X1 U2625 ( .A(n6512), .B(n6726), .C(n1384), .Y(n3785) );
  NAND2X1 U2626 ( .A(\Mem[46][27] ), .B(n6727), .Y(n1384) );
  OAI21X1 U2627 ( .A(n6507), .B(n6726), .C(n1385), .Y(n3786) );
  NAND2X1 U2628 ( .A(\Mem[46][28] ), .B(n6727), .Y(n1385) );
  OAI21X1 U2629 ( .A(n6502), .B(n6726), .C(n1386), .Y(n3787) );
  NAND2X1 U2630 ( .A(\Mem[46][29] ), .B(n6727), .Y(n1386) );
  OAI21X1 U2631 ( .A(n6492), .B(n6726), .C(n1387), .Y(n3788) );
  NAND2X1 U2632 ( .A(\Mem[46][30] ), .B(n6728), .Y(n1387) );
  OAI21X1 U2633 ( .A(n6487), .B(n6726), .C(n1388), .Y(n3789) );
  NAND2X1 U2634 ( .A(\Mem[46][31] ), .B(n6728), .Y(n1388) );
  NAND2X1 U2635 ( .A(n7010), .B(n7024), .Y(n1356) );
  OAI21X1 U2636 ( .A(n6607), .B(n6720), .C(n1390), .Y(n3790) );
  NAND2X1 U2637 ( .A(\Mem[47][0] ), .B(n6723), .Y(n1390) );
  OAI21X1 U2638 ( .A(n6552), .B(n6719), .C(n1391), .Y(n3791) );
  NAND2X1 U2639 ( .A(\Mem[47][1] ), .B(n6723), .Y(n1391) );
  OAI21X1 U2640 ( .A(n6497), .B(n6719), .C(n1392), .Y(n3792) );
  NAND2X1 U2641 ( .A(\Mem[47][2] ), .B(n6723), .Y(n1392) );
  OAI21X1 U2642 ( .A(n6482), .B(n6719), .C(n1393), .Y(n3793) );
  NAND2X1 U2643 ( .A(\Mem[47][3] ), .B(n6722), .Y(n1393) );
  OAI21X1 U2644 ( .A(n6477), .B(n6719), .C(n1394), .Y(n3794) );
  NAND2X1 U2645 ( .A(\Mem[47][4] ), .B(n6723), .Y(n1394) );
  OAI21X1 U2646 ( .A(n6472), .B(n6719), .C(n1395), .Y(n3795) );
  NAND2X1 U2647 ( .A(\Mem[47][5] ), .B(n6722), .Y(n1395) );
  OAI21X1 U2648 ( .A(n6467), .B(n6719), .C(n1396), .Y(n3796) );
  NAND2X1 U2649 ( .A(\Mem[47][6] ), .B(n6722), .Y(n1396) );
  OAI21X1 U2650 ( .A(n6462), .B(n6719), .C(n1397), .Y(n3797) );
  NAND2X1 U2651 ( .A(\Mem[47][7] ), .B(n6722), .Y(n1397) );
  OAI21X1 U2652 ( .A(n6457), .B(n6719), .C(n1398), .Y(n3798) );
  NAND2X1 U2653 ( .A(\Mem[47][8] ), .B(n6722), .Y(n1398) );
  OAI21X1 U2654 ( .A(n6452), .B(n6719), .C(n1399), .Y(n3799) );
  NAND2X1 U2655 ( .A(\Mem[47][9] ), .B(n6722), .Y(n1399) );
  OAI21X1 U2656 ( .A(n6602), .B(n6719), .C(n1400), .Y(n3800) );
  NAND2X1 U2657 ( .A(\Mem[47][10] ), .B(n6722), .Y(n1400) );
  OAI21X1 U2658 ( .A(n6597), .B(n6719), .C(n1401), .Y(n3801) );
  NAND2X1 U2659 ( .A(\Mem[47][11] ), .B(n6722), .Y(n1401) );
  OAI21X1 U2660 ( .A(n6592), .B(n6719), .C(n1402), .Y(n3802) );
  NAND2X1 U2661 ( .A(\Mem[47][12] ), .B(n6722), .Y(n1402) );
  OAI21X1 U2662 ( .A(n6587), .B(n6720), .C(n1403), .Y(n3803) );
  NAND2X1 U2663 ( .A(\Mem[47][13] ), .B(n6722), .Y(n1403) );
  OAI21X1 U2664 ( .A(n6582), .B(n6720), .C(n1404), .Y(n3804) );
  NAND2X1 U2665 ( .A(\Mem[47][14] ), .B(n6722), .Y(n1404) );
  OAI21X1 U2666 ( .A(n6577), .B(n6720), .C(n1405), .Y(n3805) );
  NAND2X1 U2667 ( .A(\Mem[47][15] ), .B(n6721), .Y(n1405) );
  OAI21X1 U2668 ( .A(n6572), .B(n6720), .C(n1406), .Y(n3806) );
  NAND2X1 U2669 ( .A(\Mem[47][16] ), .B(n6722), .Y(n1406) );
  OAI21X1 U2670 ( .A(n6567), .B(n6720), .C(n1407), .Y(n3807) );
  NAND2X1 U2671 ( .A(\Mem[47][17] ), .B(n6721), .Y(n1407) );
  OAI21X1 U2672 ( .A(n6562), .B(n6720), .C(n1408), .Y(n3808) );
  NAND2X1 U2673 ( .A(\Mem[47][18] ), .B(n6721), .Y(n1408) );
  OAI21X1 U2674 ( .A(n6557), .B(n6720), .C(n1409), .Y(n3809) );
  NAND2X1 U2675 ( .A(\Mem[47][19] ), .B(n6721), .Y(n1409) );
  OAI21X1 U2676 ( .A(n6547), .B(n6720), .C(n1410), .Y(n3810) );
  NAND2X1 U2677 ( .A(\Mem[47][20] ), .B(n6721), .Y(n1410) );
  OAI21X1 U2678 ( .A(n6542), .B(n6720), .C(n1411), .Y(n3811) );
  NAND2X1 U2679 ( .A(\Mem[47][21] ), .B(n6721), .Y(n1411) );
  OAI21X1 U2680 ( .A(n6537), .B(n6720), .C(n1412), .Y(n3812) );
  NAND2X1 U2681 ( .A(\Mem[47][22] ), .B(n6722), .Y(n1412) );
  OAI21X1 U2682 ( .A(n6532), .B(n6721), .C(n1413), .Y(n3813) );
  NAND2X1 U2683 ( .A(\Mem[47][23] ), .B(n6721), .Y(n1413) );
  OAI21X1 U2684 ( .A(n6527), .B(n6720), .C(n1414), .Y(n3814) );
  NAND2X1 U2685 ( .A(\Mem[47][24] ), .B(n6722), .Y(n1414) );
  OAI21X1 U2686 ( .A(n6522), .B(n6721), .C(n1415), .Y(n3815) );
  NAND2X1 U2687 ( .A(\Mem[47][25] ), .B(n6722), .Y(n1415) );
  OAI21X1 U2688 ( .A(n6517), .B(n6721), .C(n1416), .Y(n3816) );
  NAND2X1 U2689 ( .A(\Mem[47][26] ), .B(n6722), .Y(n1416) );
  OAI21X1 U2690 ( .A(n6512), .B(n6721), .C(n1417), .Y(n3817) );
  NAND2X1 U2691 ( .A(\Mem[47][27] ), .B(n6722), .Y(n1417) );
  OAI21X1 U2692 ( .A(n6507), .B(n6721), .C(n1418), .Y(n3818) );
  NAND2X1 U2693 ( .A(\Mem[47][28] ), .B(n6722), .Y(n1418) );
  OAI21X1 U2694 ( .A(n6502), .B(n6721), .C(n1419), .Y(n3819) );
  NAND2X1 U2695 ( .A(\Mem[47][29] ), .B(n6722), .Y(n1419) );
  OAI21X1 U2696 ( .A(n6492), .B(n6721), .C(n1420), .Y(n3820) );
  NAND2X1 U2697 ( .A(\Mem[47][30] ), .B(n6723), .Y(n1420) );
  OAI21X1 U2698 ( .A(n6487), .B(n6721), .C(n1421), .Y(n3821) );
  NAND2X1 U2699 ( .A(\Mem[47][31] ), .B(n6723), .Y(n1421) );
  NAND2X1 U2700 ( .A(n7010), .B(n7021), .Y(n1389) );
  NAND3X1 U2702 ( .A(ADDR_WR[3]), .B(n7014), .C(n80), .Y(n1422) );
  OAI21X1 U2703 ( .A(n6607), .B(n6715), .C(n1424), .Y(n3822) );
  NAND2X1 U2704 ( .A(\Mem[48][0] ), .B(n6718), .Y(n1424) );
  OAI21X1 U2705 ( .A(n6552), .B(n6714), .C(n1425), .Y(n3823) );
  NAND2X1 U2706 ( .A(\Mem[48][1] ), .B(n6718), .Y(n1425) );
  OAI21X1 U2707 ( .A(n6497), .B(n6714), .C(n1426), .Y(n3824) );
  NAND2X1 U2708 ( .A(\Mem[48][2] ), .B(n6718), .Y(n1426) );
  OAI21X1 U2709 ( .A(n6482), .B(n6714), .C(n1427), .Y(n3825) );
  NAND2X1 U2710 ( .A(\Mem[48][3] ), .B(n6717), .Y(n1427) );
  OAI21X1 U2711 ( .A(n6477), .B(n6714), .C(n1428), .Y(n3826) );
  NAND2X1 U2712 ( .A(\Mem[48][4] ), .B(n6718), .Y(n1428) );
  OAI21X1 U2713 ( .A(n6472), .B(n6714), .C(n1429), .Y(n3827) );
  NAND2X1 U2714 ( .A(\Mem[48][5] ), .B(n6717), .Y(n1429) );
  OAI21X1 U2715 ( .A(n6467), .B(n6714), .C(n1430), .Y(n3828) );
  NAND2X1 U2716 ( .A(\Mem[48][6] ), .B(n6717), .Y(n1430) );
  OAI21X1 U2717 ( .A(n6462), .B(n6714), .C(n1431), .Y(n3829) );
  NAND2X1 U2718 ( .A(\Mem[48][7] ), .B(n6717), .Y(n1431) );
  OAI21X1 U2719 ( .A(n6457), .B(n6714), .C(n1432), .Y(n3830) );
  NAND2X1 U2720 ( .A(\Mem[48][8] ), .B(n6717), .Y(n1432) );
  OAI21X1 U2721 ( .A(n6452), .B(n6714), .C(n1433), .Y(n3831) );
  NAND2X1 U2722 ( .A(\Mem[48][9] ), .B(n6717), .Y(n1433) );
  OAI21X1 U2723 ( .A(n6602), .B(n6714), .C(n1434), .Y(n3832) );
  NAND2X1 U2724 ( .A(\Mem[48][10] ), .B(n6717), .Y(n1434) );
  OAI21X1 U2725 ( .A(n6597), .B(n6714), .C(n1435), .Y(n3833) );
  NAND2X1 U2726 ( .A(\Mem[48][11] ), .B(n6717), .Y(n1435) );
  OAI21X1 U2727 ( .A(n6592), .B(n6714), .C(n1436), .Y(n3834) );
  NAND2X1 U2728 ( .A(\Mem[48][12] ), .B(n6717), .Y(n1436) );
  OAI21X1 U2729 ( .A(n6587), .B(n6715), .C(n1437), .Y(n3835) );
  NAND2X1 U2730 ( .A(\Mem[48][13] ), .B(n6717), .Y(n1437) );
  OAI21X1 U2731 ( .A(n6582), .B(n6715), .C(n1438), .Y(n3836) );
  NAND2X1 U2732 ( .A(\Mem[48][14] ), .B(n6717), .Y(n1438) );
  OAI21X1 U2733 ( .A(n6577), .B(n6715), .C(n1439), .Y(n3837) );
  NAND2X1 U2734 ( .A(\Mem[48][15] ), .B(n6716), .Y(n1439) );
  OAI21X1 U2735 ( .A(n6572), .B(n6715), .C(n1440), .Y(n3838) );
  NAND2X1 U2736 ( .A(\Mem[48][16] ), .B(n6717), .Y(n1440) );
  OAI21X1 U2737 ( .A(n6567), .B(n6715), .C(n1441), .Y(n3839) );
  NAND2X1 U2738 ( .A(\Mem[48][17] ), .B(n6716), .Y(n1441) );
  OAI21X1 U2739 ( .A(n6562), .B(n6715), .C(n1442), .Y(n3840) );
  NAND2X1 U2740 ( .A(\Mem[48][18] ), .B(n6716), .Y(n1442) );
  OAI21X1 U2741 ( .A(n6557), .B(n6715), .C(n1443), .Y(n3841) );
  NAND2X1 U2742 ( .A(\Mem[48][19] ), .B(n6716), .Y(n1443) );
  OAI21X1 U2743 ( .A(n6547), .B(n6715), .C(n1444), .Y(n3842) );
  NAND2X1 U2744 ( .A(\Mem[48][20] ), .B(n6716), .Y(n1444) );
  OAI21X1 U2745 ( .A(n6542), .B(n6715), .C(n1445), .Y(n3843) );
  NAND2X1 U2746 ( .A(\Mem[48][21] ), .B(n6716), .Y(n1445) );
  OAI21X1 U2747 ( .A(n6537), .B(n6715), .C(n1446), .Y(n3844) );
  NAND2X1 U2748 ( .A(\Mem[48][22] ), .B(n6717), .Y(n1446) );
  OAI21X1 U2749 ( .A(n6532), .B(n6716), .C(n1447), .Y(n3845) );
  NAND2X1 U2750 ( .A(\Mem[48][23] ), .B(n6716), .Y(n1447) );
  OAI21X1 U2751 ( .A(n6527), .B(n6715), .C(n1448), .Y(n3846) );
  NAND2X1 U2752 ( .A(\Mem[48][24] ), .B(n6717), .Y(n1448) );
  OAI21X1 U2753 ( .A(n6522), .B(n6716), .C(n1449), .Y(n3847) );
  NAND2X1 U2754 ( .A(\Mem[48][25] ), .B(n6717), .Y(n1449) );
  OAI21X1 U2755 ( .A(n6517), .B(n6716), .C(n1450), .Y(n3848) );
  NAND2X1 U2756 ( .A(\Mem[48][26] ), .B(n6717), .Y(n1450) );
  OAI21X1 U2757 ( .A(n6512), .B(n6716), .C(n1451), .Y(n3849) );
  NAND2X1 U2758 ( .A(\Mem[48][27] ), .B(n6717), .Y(n1451) );
  OAI21X1 U2759 ( .A(n6507), .B(n6716), .C(n1452), .Y(n3850) );
  NAND2X1 U2760 ( .A(\Mem[48][28] ), .B(n6717), .Y(n1452) );
  OAI21X1 U2761 ( .A(n6502), .B(n6716), .C(n1453), .Y(n3851) );
  NAND2X1 U2762 ( .A(\Mem[48][29] ), .B(n6717), .Y(n1453) );
  OAI21X1 U2763 ( .A(n6492), .B(n6716), .C(n1454), .Y(n3852) );
  NAND2X1 U2764 ( .A(\Mem[48][30] ), .B(n6718), .Y(n1454) );
  OAI21X1 U2765 ( .A(n6487), .B(n6716), .C(n1455), .Y(n3853) );
  NAND2X1 U2766 ( .A(\Mem[48][31] ), .B(n6718), .Y(n1455) );
  NAND2X1 U2767 ( .A(n7009), .B(n7016), .Y(n1423) );
  OAI21X1 U2768 ( .A(n6607), .B(n6710), .C(n1458), .Y(n3854) );
  NAND2X1 U2769 ( .A(\Mem[49][0] ), .B(n6713), .Y(n1458) );
  OAI21X1 U2770 ( .A(n6552), .B(n6709), .C(n1459), .Y(n3855) );
  NAND2X1 U2771 ( .A(\Mem[49][1] ), .B(n6713), .Y(n1459) );
  OAI21X1 U2772 ( .A(n6497), .B(n6709), .C(n1460), .Y(n3856) );
  NAND2X1 U2773 ( .A(\Mem[49][2] ), .B(n6713), .Y(n1460) );
  OAI21X1 U2774 ( .A(n6482), .B(n6709), .C(n1461), .Y(n3857) );
  NAND2X1 U2775 ( .A(\Mem[49][3] ), .B(n6712), .Y(n1461) );
  OAI21X1 U2776 ( .A(n6477), .B(n6709), .C(n1462), .Y(n3858) );
  NAND2X1 U2777 ( .A(\Mem[49][4] ), .B(n6713), .Y(n1462) );
  OAI21X1 U2778 ( .A(n6472), .B(n6709), .C(n1463), .Y(n3859) );
  NAND2X1 U2779 ( .A(\Mem[49][5] ), .B(n6712), .Y(n1463) );
  OAI21X1 U2780 ( .A(n6467), .B(n6709), .C(n1464), .Y(n3860) );
  NAND2X1 U2781 ( .A(\Mem[49][6] ), .B(n6712), .Y(n1464) );
  OAI21X1 U2782 ( .A(n6462), .B(n6709), .C(n1465), .Y(n3861) );
  NAND2X1 U2783 ( .A(\Mem[49][7] ), .B(n6712), .Y(n1465) );
  OAI21X1 U2784 ( .A(n6457), .B(n6709), .C(n1466), .Y(n3862) );
  NAND2X1 U2785 ( .A(\Mem[49][8] ), .B(n6712), .Y(n1466) );
  OAI21X1 U2786 ( .A(n6452), .B(n6709), .C(n1467), .Y(n3863) );
  NAND2X1 U2787 ( .A(\Mem[49][9] ), .B(n6712), .Y(n1467) );
  OAI21X1 U2788 ( .A(n6602), .B(n6709), .C(n1468), .Y(n3864) );
  NAND2X1 U2789 ( .A(\Mem[49][10] ), .B(n6712), .Y(n1468) );
  OAI21X1 U2790 ( .A(n6597), .B(n6709), .C(n1469), .Y(n3865) );
  NAND2X1 U2791 ( .A(\Mem[49][11] ), .B(n6712), .Y(n1469) );
  OAI21X1 U2792 ( .A(n6592), .B(n6709), .C(n1470), .Y(n3866) );
  NAND2X1 U2793 ( .A(\Mem[49][12] ), .B(n6712), .Y(n1470) );
  OAI21X1 U2794 ( .A(n6587), .B(n6710), .C(n1471), .Y(n3867) );
  NAND2X1 U2795 ( .A(\Mem[49][13] ), .B(n6712), .Y(n1471) );
  OAI21X1 U2796 ( .A(n6582), .B(n6710), .C(n1472), .Y(n3868) );
  NAND2X1 U2797 ( .A(\Mem[49][14] ), .B(n6712), .Y(n1472) );
  OAI21X1 U2798 ( .A(n6577), .B(n6710), .C(n1473), .Y(n3869) );
  NAND2X1 U2799 ( .A(\Mem[49][15] ), .B(n6711), .Y(n1473) );
  OAI21X1 U2800 ( .A(n6572), .B(n6710), .C(n1474), .Y(n3870) );
  NAND2X1 U2801 ( .A(\Mem[49][16] ), .B(n6712), .Y(n1474) );
  OAI21X1 U2802 ( .A(n6567), .B(n6710), .C(n1475), .Y(n3871) );
  NAND2X1 U2803 ( .A(\Mem[49][17] ), .B(n6711), .Y(n1475) );
  OAI21X1 U2804 ( .A(n6562), .B(n6710), .C(n1476), .Y(n3872) );
  NAND2X1 U2805 ( .A(\Mem[49][18] ), .B(n6711), .Y(n1476) );
  OAI21X1 U2806 ( .A(n6557), .B(n6710), .C(n1477), .Y(n3873) );
  NAND2X1 U2807 ( .A(\Mem[49][19] ), .B(n6711), .Y(n1477) );
  OAI21X1 U2808 ( .A(n6547), .B(n6710), .C(n1478), .Y(n3874) );
  NAND2X1 U2809 ( .A(\Mem[49][20] ), .B(n6711), .Y(n1478) );
  OAI21X1 U2810 ( .A(n6542), .B(n6710), .C(n1479), .Y(n3875) );
  NAND2X1 U2811 ( .A(\Mem[49][21] ), .B(n6711), .Y(n1479) );
  OAI21X1 U2812 ( .A(n6537), .B(n6710), .C(n1480), .Y(n3876) );
  NAND2X1 U2813 ( .A(\Mem[49][22] ), .B(n6712), .Y(n1480) );
  OAI21X1 U2814 ( .A(n6532), .B(n6711), .C(n1481), .Y(n3877) );
  NAND2X1 U2815 ( .A(\Mem[49][23] ), .B(n6711), .Y(n1481) );
  OAI21X1 U2816 ( .A(n6527), .B(n6710), .C(n1482), .Y(n3878) );
  NAND2X1 U2817 ( .A(\Mem[49][24] ), .B(n6712), .Y(n1482) );
  OAI21X1 U2818 ( .A(n6522), .B(n6711), .C(n1483), .Y(n3879) );
  NAND2X1 U2819 ( .A(\Mem[49][25] ), .B(n6712), .Y(n1483) );
  OAI21X1 U2820 ( .A(n6517), .B(n6711), .C(n1484), .Y(n3880) );
  NAND2X1 U2821 ( .A(\Mem[49][26] ), .B(n6712), .Y(n1484) );
  OAI21X1 U2822 ( .A(n6512), .B(n6711), .C(n1485), .Y(n3881) );
  NAND2X1 U2823 ( .A(\Mem[49][27] ), .B(n6712), .Y(n1485) );
  OAI21X1 U2824 ( .A(n6507), .B(n6711), .C(n1486), .Y(n3882) );
  NAND2X1 U2825 ( .A(\Mem[49][28] ), .B(n6712), .Y(n1486) );
  OAI21X1 U2826 ( .A(n6502), .B(n6711), .C(n1487), .Y(n3883) );
  NAND2X1 U2827 ( .A(\Mem[49][29] ), .B(n6712), .Y(n1487) );
  OAI21X1 U2828 ( .A(n6492), .B(n6711), .C(n1488), .Y(n3884) );
  NAND2X1 U2829 ( .A(\Mem[49][30] ), .B(n6713), .Y(n1488) );
  OAI21X1 U2830 ( .A(n6487), .B(n6711), .C(n1489), .Y(n3885) );
  NAND2X1 U2831 ( .A(\Mem[49][31] ), .B(n6713), .Y(n1489) );
  NAND2X1 U2832 ( .A(n7009), .B(n7017), .Y(n1457) );
  OAI21X1 U2833 ( .A(n6607), .B(n6705), .C(n1491), .Y(n3886) );
  NAND2X1 U2834 ( .A(\Mem[50][0] ), .B(n6708), .Y(n1491) );
  OAI21X1 U2835 ( .A(n6552), .B(n6704), .C(n1492), .Y(n3887) );
  NAND2X1 U2836 ( .A(\Mem[50][1] ), .B(n6708), .Y(n1492) );
  OAI21X1 U2837 ( .A(n6497), .B(n6704), .C(n1493), .Y(n3888) );
  NAND2X1 U2838 ( .A(\Mem[50][2] ), .B(n6708), .Y(n1493) );
  OAI21X1 U2839 ( .A(n6482), .B(n6704), .C(n1494), .Y(n3889) );
  NAND2X1 U2840 ( .A(\Mem[50][3] ), .B(n6707), .Y(n1494) );
  OAI21X1 U2841 ( .A(n6477), .B(n6704), .C(n1495), .Y(n3890) );
  NAND2X1 U2842 ( .A(\Mem[50][4] ), .B(n6708), .Y(n1495) );
  OAI21X1 U2843 ( .A(n6472), .B(n6704), .C(n1496), .Y(n3891) );
  NAND2X1 U2844 ( .A(\Mem[50][5] ), .B(n6707), .Y(n1496) );
  OAI21X1 U2845 ( .A(n6467), .B(n6704), .C(n1497), .Y(n3892) );
  NAND2X1 U2846 ( .A(\Mem[50][6] ), .B(n6707), .Y(n1497) );
  OAI21X1 U2847 ( .A(n6462), .B(n6704), .C(n1498), .Y(n3893) );
  NAND2X1 U2848 ( .A(\Mem[50][7] ), .B(n6707), .Y(n1498) );
  OAI21X1 U2849 ( .A(n6457), .B(n6704), .C(n1499), .Y(n3894) );
  NAND2X1 U2850 ( .A(\Mem[50][8] ), .B(n6707), .Y(n1499) );
  OAI21X1 U2851 ( .A(n6452), .B(n6704), .C(n1500), .Y(n3895) );
  NAND2X1 U2852 ( .A(\Mem[50][9] ), .B(n6707), .Y(n1500) );
  OAI21X1 U2853 ( .A(n6602), .B(n6704), .C(n1501), .Y(n3896) );
  NAND2X1 U2854 ( .A(\Mem[50][10] ), .B(n6707), .Y(n1501) );
  OAI21X1 U2855 ( .A(n6597), .B(n6704), .C(n1502), .Y(n3897) );
  NAND2X1 U2856 ( .A(\Mem[50][11] ), .B(n6707), .Y(n1502) );
  OAI21X1 U2857 ( .A(n6592), .B(n6704), .C(n1503), .Y(n3898) );
  NAND2X1 U2858 ( .A(\Mem[50][12] ), .B(n6707), .Y(n1503) );
  OAI21X1 U2859 ( .A(n6587), .B(n6705), .C(n1504), .Y(n3899) );
  NAND2X1 U2860 ( .A(\Mem[50][13] ), .B(n6707), .Y(n1504) );
  OAI21X1 U2861 ( .A(n6582), .B(n6705), .C(n1505), .Y(n3900) );
  NAND2X1 U2862 ( .A(\Mem[50][14] ), .B(n6707), .Y(n1505) );
  OAI21X1 U2863 ( .A(n6577), .B(n6705), .C(n1506), .Y(n3901) );
  NAND2X1 U2864 ( .A(\Mem[50][15] ), .B(n6706), .Y(n1506) );
  OAI21X1 U2865 ( .A(n6572), .B(n6705), .C(n1507), .Y(n3902) );
  NAND2X1 U2866 ( .A(\Mem[50][16] ), .B(n6707), .Y(n1507) );
  OAI21X1 U2867 ( .A(n6567), .B(n6705), .C(n1508), .Y(n3903) );
  NAND2X1 U2868 ( .A(\Mem[50][17] ), .B(n6706), .Y(n1508) );
  OAI21X1 U2869 ( .A(n6562), .B(n6705), .C(n1509), .Y(n3904) );
  NAND2X1 U2870 ( .A(\Mem[50][18] ), .B(n6706), .Y(n1509) );
  OAI21X1 U2871 ( .A(n6557), .B(n6705), .C(n1510), .Y(n3905) );
  NAND2X1 U2872 ( .A(\Mem[50][19] ), .B(n6706), .Y(n1510) );
  OAI21X1 U2873 ( .A(n6547), .B(n6705), .C(n1511), .Y(n3906) );
  NAND2X1 U2874 ( .A(\Mem[50][20] ), .B(n6706), .Y(n1511) );
  OAI21X1 U2875 ( .A(n6542), .B(n6705), .C(n1512), .Y(n3907) );
  NAND2X1 U2876 ( .A(\Mem[50][21] ), .B(n6706), .Y(n1512) );
  OAI21X1 U2877 ( .A(n6537), .B(n6705), .C(n1513), .Y(n3908) );
  NAND2X1 U2878 ( .A(\Mem[50][22] ), .B(n6707), .Y(n1513) );
  OAI21X1 U2879 ( .A(n6532), .B(n6706), .C(n1514), .Y(n3909) );
  NAND2X1 U2880 ( .A(\Mem[50][23] ), .B(n6706), .Y(n1514) );
  OAI21X1 U2881 ( .A(n6527), .B(n6705), .C(n1515), .Y(n3910) );
  NAND2X1 U2882 ( .A(\Mem[50][24] ), .B(n6707), .Y(n1515) );
  OAI21X1 U2883 ( .A(n6522), .B(n6706), .C(n1516), .Y(n3911) );
  NAND2X1 U2884 ( .A(\Mem[50][25] ), .B(n6707), .Y(n1516) );
  OAI21X1 U2885 ( .A(n6517), .B(n6706), .C(n1517), .Y(n3912) );
  NAND2X1 U2886 ( .A(\Mem[50][26] ), .B(n6707), .Y(n1517) );
  OAI21X1 U2887 ( .A(n6512), .B(n6706), .C(n1518), .Y(n3913) );
  NAND2X1 U2888 ( .A(\Mem[50][27] ), .B(n6707), .Y(n1518) );
  OAI21X1 U2889 ( .A(n6507), .B(n6706), .C(n1519), .Y(n3914) );
  NAND2X1 U2890 ( .A(\Mem[50][28] ), .B(n6707), .Y(n1519) );
  OAI21X1 U2891 ( .A(n6502), .B(n6706), .C(n1520), .Y(n3915) );
  NAND2X1 U2892 ( .A(\Mem[50][29] ), .B(n6707), .Y(n1520) );
  OAI21X1 U2893 ( .A(n6492), .B(n6706), .C(n1521), .Y(n3916) );
  NAND2X1 U2894 ( .A(\Mem[50][30] ), .B(n6708), .Y(n1521) );
  OAI21X1 U2895 ( .A(n6487), .B(n6706), .C(n1522), .Y(n3917) );
  NAND2X1 U2896 ( .A(\Mem[50][31] ), .B(n6708), .Y(n1522) );
  NAND2X1 U2897 ( .A(n7009), .B(n7018), .Y(n1490) );
  OAI21X1 U2898 ( .A(n6607), .B(n6700), .C(n1524), .Y(n3918) );
  NAND2X1 U2899 ( .A(\Mem[51][0] ), .B(n6703), .Y(n1524) );
  OAI21X1 U2900 ( .A(n6552), .B(n6699), .C(n1525), .Y(n3919) );
  NAND2X1 U2901 ( .A(\Mem[51][1] ), .B(n6703), .Y(n1525) );
  OAI21X1 U2902 ( .A(n6497), .B(n6699), .C(n1526), .Y(n3920) );
  NAND2X1 U2903 ( .A(\Mem[51][2] ), .B(n6703), .Y(n1526) );
  OAI21X1 U2904 ( .A(n6482), .B(n6699), .C(n1527), .Y(n3921) );
  NAND2X1 U2905 ( .A(\Mem[51][3] ), .B(n6702), .Y(n1527) );
  OAI21X1 U2906 ( .A(n6477), .B(n6699), .C(n1528), .Y(n3922) );
  NAND2X1 U2907 ( .A(\Mem[51][4] ), .B(n6703), .Y(n1528) );
  OAI21X1 U2908 ( .A(n6472), .B(n6699), .C(n1529), .Y(n3923) );
  NAND2X1 U2909 ( .A(\Mem[51][5] ), .B(n6702), .Y(n1529) );
  OAI21X1 U2910 ( .A(n6467), .B(n6699), .C(n1530), .Y(n3924) );
  NAND2X1 U2911 ( .A(\Mem[51][6] ), .B(n6702), .Y(n1530) );
  OAI21X1 U2912 ( .A(n6462), .B(n6699), .C(n1531), .Y(n3925) );
  NAND2X1 U2913 ( .A(\Mem[51][7] ), .B(n6702), .Y(n1531) );
  OAI21X1 U2914 ( .A(n6457), .B(n6699), .C(n1532), .Y(n3926) );
  NAND2X1 U2915 ( .A(\Mem[51][8] ), .B(n6702), .Y(n1532) );
  OAI21X1 U2916 ( .A(n6452), .B(n6699), .C(n1533), .Y(n3927) );
  NAND2X1 U2917 ( .A(\Mem[51][9] ), .B(n6702), .Y(n1533) );
  OAI21X1 U2918 ( .A(n6602), .B(n6699), .C(n1534), .Y(n3928) );
  NAND2X1 U2919 ( .A(\Mem[51][10] ), .B(n6702), .Y(n1534) );
  OAI21X1 U2920 ( .A(n6597), .B(n6699), .C(n1535), .Y(n3929) );
  NAND2X1 U2921 ( .A(\Mem[51][11] ), .B(n6702), .Y(n1535) );
  OAI21X1 U2922 ( .A(n6592), .B(n6699), .C(n1536), .Y(n3930) );
  NAND2X1 U2923 ( .A(\Mem[51][12] ), .B(n6702), .Y(n1536) );
  OAI21X1 U2924 ( .A(n6587), .B(n6700), .C(n1537), .Y(n3931) );
  NAND2X1 U2925 ( .A(\Mem[51][13] ), .B(n6702), .Y(n1537) );
  OAI21X1 U2926 ( .A(n6582), .B(n6700), .C(n1538), .Y(n3932) );
  NAND2X1 U2927 ( .A(\Mem[51][14] ), .B(n6702), .Y(n1538) );
  OAI21X1 U2928 ( .A(n6577), .B(n6700), .C(n1539), .Y(n3933) );
  NAND2X1 U2929 ( .A(\Mem[51][15] ), .B(n6701), .Y(n1539) );
  OAI21X1 U2930 ( .A(n6572), .B(n6700), .C(n1540), .Y(n3934) );
  NAND2X1 U2931 ( .A(\Mem[51][16] ), .B(n6702), .Y(n1540) );
  OAI21X1 U2932 ( .A(n6567), .B(n6700), .C(n1541), .Y(n3935) );
  NAND2X1 U2933 ( .A(\Mem[51][17] ), .B(n6701), .Y(n1541) );
  OAI21X1 U2934 ( .A(n6562), .B(n6700), .C(n1542), .Y(n3936) );
  NAND2X1 U2935 ( .A(\Mem[51][18] ), .B(n6701), .Y(n1542) );
  OAI21X1 U2936 ( .A(n6557), .B(n6700), .C(n1543), .Y(n3937) );
  NAND2X1 U2937 ( .A(\Mem[51][19] ), .B(n6701), .Y(n1543) );
  OAI21X1 U2938 ( .A(n6547), .B(n6700), .C(n1544), .Y(n3938) );
  NAND2X1 U2939 ( .A(\Mem[51][20] ), .B(n6701), .Y(n1544) );
  OAI21X1 U2940 ( .A(n6542), .B(n6700), .C(n1545), .Y(n3939) );
  NAND2X1 U2941 ( .A(\Mem[51][21] ), .B(n6701), .Y(n1545) );
  OAI21X1 U2942 ( .A(n6537), .B(n6700), .C(n1546), .Y(n3940) );
  NAND2X1 U2943 ( .A(\Mem[51][22] ), .B(n6702), .Y(n1546) );
  OAI21X1 U2944 ( .A(n6532), .B(n6701), .C(n1547), .Y(n3941) );
  NAND2X1 U2945 ( .A(\Mem[51][23] ), .B(n6701), .Y(n1547) );
  OAI21X1 U2946 ( .A(n6527), .B(n6700), .C(n1548), .Y(n3942) );
  NAND2X1 U2947 ( .A(\Mem[51][24] ), .B(n6702), .Y(n1548) );
  OAI21X1 U2948 ( .A(n6522), .B(n6701), .C(n1549), .Y(n3943) );
  NAND2X1 U2949 ( .A(\Mem[51][25] ), .B(n6702), .Y(n1549) );
  OAI21X1 U2950 ( .A(n6517), .B(n6701), .C(n1550), .Y(n3944) );
  NAND2X1 U2951 ( .A(\Mem[51][26] ), .B(n6702), .Y(n1550) );
  OAI21X1 U2952 ( .A(n6512), .B(n6701), .C(n1551), .Y(n3945) );
  NAND2X1 U2953 ( .A(\Mem[51][27] ), .B(n6702), .Y(n1551) );
  OAI21X1 U2954 ( .A(n6507), .B(n6701), .C(n1552), .Y(n3946) );
  NAND2X1 U2955 ( .A(\Mem[51][28] ), .B(n6702), .Y(n1552) );
  OAI21X1 U2956 ( .A(n6502), .B(n6701), .C(n1553), .Y(n3947) );
  NAND2X1 U2957 ( .A(\Mem[51][29] ), .B(n6702), .Y(n1553) );
  OAI21X1 U2958 ( .A(n6492), .B(n6701), .C(n1554), .Y(n3948) );
  NAND2X1 U2959 ( .A(\Mem[51][30] ), .B(n6703), .Y(n1554) );
  OAI21X1 U2960 ( .A(n6487), .B(n6701), .C(n1555), .Y(n3949) );
  NAND2X1 U2961 ( .A(\Mem[51][31] ), .B(n6703), .Y(n1555) );
  NAND2X1 U2962 ( .A(n7009), .B(n7019), .Y(n1523) );
  OAI21X1 U2963 ( .A(n6607), .B(n6695), .C(n1557), .Y(n3950) );
  NAND2X1 U2964 ( .A(\Mem[52][0] ), .B(n6698), .Y(n1557) );
  OAI21X1 U2965 ( .A(n6552), .B(n6694), .C(n1558), .Y(n3951) );
  NAND2X1 U2966 ( .A(\Mem[52][1] ), .B(n6698), .Y(n1558) );
  OAI21X1 U2967 ( .A(n6497), .B(n6694), .C(n1559), .Y(n3952) );
  NAND2X1 U2968 ( .A(\Mem[52][2] ), .B(n6698), .Y(n1559) );
  OAI21X1 U2969 ( .A(n6482), .B(n6694), .C(n1560), .Y(n3953) );
  NAND2X1 U2970 ( .A(\Mem[52][3] ), .B(n6697), .Y(n1560) );
  OAI21X1 U2971 ( .A(n6477), .B(n6694), .C(n1561), .Y(n3954) );
  NAND2X1 U2972 ( .A(\Mem[52][4] ), .B(n6698), .Y(n1561) );
  OAI21X1 U2973 ( .A(n6472), .B(n6694), .C(n1562), .Y(n3955) );
  NAND2X1 U2974 ( .A(\Mem[52][5] ), .B(n6697), .Y(n1562) );
  OAI21X1 U2975 ( .A(n6467), .B(n6694), .C(n1563), .Y(n3956) );
  NAND2X1 U2976 ( .A(\Mem[52][6] ), .B(n6697), .Y(n1563) );
  OAI21X1 U2977 ( .A(n6462), .B(n6694), .C(n1564), .Y(n3957) );
  NAND2X1 U2978 ( .A(\Mem[52][7] ), .B(n6697), .Y(n1564) );
  OAI21X1 U2979 ( .A(n6457), .B(n6694), .C(n1565), .Y(n3958) );
  NAND2X1 U2980 ( .A(\Mem[52][8] ), .B(n6697), .Y(n1565) );
  OAI21X1 U2981 ( .A(n6452), .B(n6694), .C(n1566), .Y(n3959) );
  NAND2X1 U2982 ( .A(\Mem[52][9] ), .B(n6697), .Y(n1566) );
  OAI21X1 U2983 ( .A(n6602), .B(n6694), .C(n1567), .Y(n3960) );
  NAND2X1 U2984 ( .A(\Mem[52][10] ), .B(n6697), .Y(n1567) );
  OAI21X1 U2985 ( .A(n6597), .B(n6694), .C(n1568), .Y(n3961) );
  NAND2X1 U2986 ( .A(\Mem[52][11] ), .B(n6697), .Y(n1568) );
  OAI21X1 U2987 ( .A(n6592), .B(n6694), .C(n1569), .Y(n3962) );
  NAND2X1 U2988 ( .A(\Mem[52][12] ), .B(n6697), .Y(n1569) );
  OAI21X1 U2989 ( .A(n6587), .B(n6695), .C(n1570), .Y(n3963) );
  NAND2X1 U2990 ( .A(\Mem[52][13] ), .B(n6697), .Y(n1570) );
  OAI21X1 U2991 ( .A(n6582), .B(n6695), .C(n1571), .Y(n3964) );
  NAND2X1 U2992 ( .A(\Mem[52][14] ), .B(n6697), .Y(n1571) );
  OAI21X1 U2993 ( .A(n6577), .B(n6695), .C(n1572), .Y(n3965) );
  NAND2X1 U2994 ( .A(\Mem[52][15] ), .B(n6696), .Y(n1572) );
  OAI21X1 U2995 ( .A(n6572), .B(n6695), .C(n1573), .Y(n3966) );
  NAND2X1 U2996 ( .A(\Mem[52][16] ), .B(n6697), .Y(n1573) );
  OAI21X1 U2997 ( .A(n6567), .B(n6695), .C(n1574), .Y(n3967) );
  NAND2X1 U2998 ( .A(\Mem[52][17] ), .B(n6696), .Y(n1574) );
  OAI21X1 U2999 ( .A(n6562), .B(n6695), .C(n1575), .Y(n3968) );
  NAND2X1 U3000 ( .A(\Mem[52][18] ), .B(n6696), .Y(n1575) );
  OAI21X1 U3001 ( .A(n6557), .B(n6695), .C(n1576), .Y(n3969) );
  NAND2X1 U3002 ( .A(\Mem[52][19] ), .B(n6696), .Y(n1576) );
  OAI21X1 U3003 ( .A(n6547), .B(n6695), .C(n1577), .Y(n3970) );
  NAND2X1 U3004 ( .A(\Mem[52][20] ), .B(n6696), .Y(n1577) );
  OAI21X1 U3005 ( .A(n6542), .B(n6695), .C(n1578), .Y(n3971) );
  NAND2X1 U3006 ( .A(\Mem[52][21] ), .B(n6696), .Y(n1578) );
  OAI21X1 U3007 ( .A(n6537), .B(n6695), .C(n1579), .Y(n3972) );
  NAND2X1 U3008 ( .A(\Mem[52][22] ), .B(n6697), .Y(n1579) );
  OAI21X1 U3009 ( .A(n6532), .B(n6696), .C(n1580), .Y(n3973) );
  NAND2X1 U3010 ( .A(\Mem[52][23] ), .B(n6696), .Y(n1580) );
  OAI21X1 U3011 ( .A(n6527), .B(n6695), .C(n1581), .Y(n3974) );
  NAND2X1 U3012 ( .A(\Mem[52][24] ), .B(n6697), .Y(n1581) );
  OAI21X1 U3013 ( .A(n6522), .B(n6696), .C(n1582), .Y(n3975) );
  NAND2X1 U3014 ( .A(\Mem[52][25] ), .B(n6697), .Y(n1582) );
  OAI21X1 U3015 ( .A(n6517), .B(n6696), .C(n1583), .Y(n3976) );
  NAND2X1 U3016 ( .A(\Mem[52][26] ), .B(n6697), .Y(n1583) );
  OAI21X1 U3017 ( .A(n6512), .B(n6696), .C(n1584), .Y(n3977) );
  NAND2X1 U3018 ( .A(\Mem[52][27] ), .B(n6697), .Y(n1584) );
  OAI21X1 U3019 ( .A(n6507), .B(n6696), .C(n1585), .Y(n3978) );
  NAND2X1 U3020 ( .A(\Mem[52][28] ), .B(n6697), .Y(n1585) );
  OAI21X1 U3021 ( .A(n6502), .B(n6696), .C(n1586), .Y(n3979) );
  NAND2X1 U3022 ( .A(\Mem[52][29] ), .B(n6697), .Y(n1586) );
  OAI21X1 U3023 ( .A(n6492), .B(n6696), .C(n1587), .Y(n3980) );
  NAND2X1 U3024 ( .A(\Mem[52][30] ), .B(n6698), .Y(n1587) );
  OAI21X1 U3025 ( .A(n6487), .B(n6696), .C(n1588), .Y(n3981) );
  NAND2X1 U3026 ( .A(\Mem[52][31] ), .B(n6698), .Y(n1588) );
  NAND2X1 U3027 ( .A(n7009), .B(n7022), .Y(n1556) );
  OAI21X1 U3028 ( .A(n6607), .B(n6690), .C(n1590), .Y(n3982) );
  NAND2X1 U3029 ( .A(\Mem[53][0] ), .B(n6693), .Y(n1590) );
  OAI21X1 U3030 ( .A(n6552), .B(n6689), .C(n1591), .Y(n3983) );
  NAND2X1 U3031 ( .A(\Mem[53][1] ), .B(n6693), .Y(n1591) );
  OAI21X1 U3032 ( .A(n6497), .B(n6689), .C(n1592), .Y(n3984) );
  NAND2X1 U3033 ( .A(\Mem[53][2] ), .B(n6693), .Y(n1592) );
  OAI21X1 U3034 ( .A(n6482), .B(n6689), .C(n1593), .Y(n3985) );
  NAND2X1 U3035 ( .A(\Mem[53][3] ), .B(n6692), .Y(n1593) );
  OAI21X1 U3036 ( .A(n6477), .B(n6689), .C(n1594), .Y(n3986) );
  NAND2X1 U3037 ( .A(\Mem[53][4] ), .B(n6693), .Y(n1594) );
  OAI21X1 U3038 ( .A(n6472), .B(n6689), .C(n1595), .Y(n3987) );
  NAND2X1 U3039 ( .A(\Mem[53][5] ), .B(n6692), .Y(n1595) );
  OAI21X1 U3040 ( .A(n6467), .B(n6689), .C(n1596), .Y(n3988) );
  NAND2X1 U3041 ( .A(\Mem[53][6] ), .B(n6692), .Y(n1596) );
  OAI21X1 U3042 ( .A(n6462), .B(n6689), .C(n1597), .Y(n3989) );
  NAND2X1 U3043 ( .A(\Mem[53][7] ), .B(n6692), .Y(n1597) );
  OAI21X1 U3044 ( .A(n6457), .B(n6689), .C(n1598), .Y(n3990) );
  NAND2X1 U3045 ( .A(\Mem[53][8] ), .B(n6692), .Y(n1598) );
  OAI21X1 U3046 ( .A(n6452), .B(n6689), .C(n1599), .Y(n3991) );
  NAND2X1 U3047 ( .A(\Mem[53][9] ), .B(n6692), .Y(n1599) );
  OAI21X1 U3048 ( .A(n6602), .B(n6689), .C(n1600), .Y(n3992) );
  NAND2X1 U3049 ( .A(\Mem[53][10] ), .B(n6692), .Y(n1600) );
  OAI21X1 U3050 ( .A(n6597), .B(n6689), .C(n1601), .Y(n3993) );
  NAND2X1 U3051 ( .A(\Mem[53][11] ), .B(n6692), .Y(n1601) );
  OAI21X1 U3052 ( .A(n6592), .B(n6689), .C(n1602), .Y(n3994) );
  NAND2X1 U3053 ( .A(\Mem[53][12] ), .B(n6692), .Y(n1602) );
  OAI21X1 U3054 ( .A(n6587), .B(n6690), .C(n1603), .Y(n3995) );
  NAND2X1 U3055 ( .A(\Mem[53][13] ), .B(n6692), .Y(n1603) );
  OAI21X1 U3056 ( .A(n6582), .B(n6690), .C(n1604), .Y(n3996) );
  NAND2X1 U3057 ( .A(\Mem[53][14] ), .B(n6692), .Y(n1604) );
  OAI21X1 U3058 ( .A(n6577), .B(n6690), .C(n1605), .Y(n3997) );
  NAND2X1 U3059 ( .A(\Mem[53][15] ), .B(n6691), .Y(n1605) );
  OAI21X1 U3060 ( .A(n6572), .B(n6690), .C(n1606), .Y(n3998) );
  NAND2X1 U3061 ( .A(\Mem[53][16] ), .B(n6692), .Y(n1606) );
  OAI21X1 U3062 ( .A(n6567), .B(n6690), .C(n1607), .Y(n3999) );
  NAND2X1 U3063 ( .A(\Mem[53][17] ), .B(n6691), .Y(n1607) );
  OAI21X1 U3064 ( .A(n6562), .B(n6690), .C(n1608), .Y(n4000) );
  NAND2X1 U3065 ( .A(\Mem[53][18] ), .B(n6691), .Y(n1608) );
  OAI21X1 U3066 ( .A(n6557), .B(n6690), .C(n1609), .Y(n4001) );
  NAND2X1 U3067 ( .A(\Mem[53][19] ), .B(n6691), .Y(n1609) );
  OAI21X1 U3068 ( .A(n6547), .B(n6690), .C(n1610), .Y(n4002) );
  NAND2X1 U3069 ( .A(\Mem[53][20] ), .B(n6691), .Y(n1610) );
  OAI21X1 U3070 ( .A(n6542), .B(n6690), .C(n1611), .Y(n4003) );
  NAND2X1 U3071 ( .A(\Mem[53][21] ), .B(n6691), .Y(n1611) );
  OAI21X1 U3072 ( .A(n6537), .B(n6690), .C(n1612), .Y(n4004) );
  NAND2X1 U3073 ( .A(\Mem[53][22] ), .B(n6692), .Y(n1612) );
  OAI21X1 U3074 ( .A(n6532), .B(n6691), .C(n1613), .Y(n4005) );
  NAND2X1 U3075 ( .A(\Mem[53][23] ), .B(n6691), .Y(n1613) );
  OAI21X1 U3076 ( .A(n6527), .B(n6690), .C(n1614), .Y(n4006) );
  NAND2X1 U3077 ( .A(\Mem[53][24] ), .B(n6692), .Y(n1614) );
  OAI21X1 U3078 ( .A(n6522), .B(n6691), .C(n1615), .Y(n4007) );
  NAND2X1 U3079 ( .A(\Mem[53][25] ), .B(n6692), .Y(n1615) );
  OAI21X1 U3080 ( .A(n6517), .B(n6691), .C(n1616), .Y(n4008) );
  NAND2X1 U3081 ( .A(\Mem[53][26] ), .B(n6692), .Y(n1616) );
  OAI21X1 U3082 ( .A(n6512), .B(n6691), .C(n1617), .Y(n4009) );
  NAND2X1 U3083 ( .A(\Mem[53][27] ), .B(n6692), .Y(n1617) );
  OAI21X1 U3084 ( .A(n6507), .B(n6691), .C(n1618), .Y(n4010) );
  NAND2X1 U3085 ( .A(\Mem[53][28] ), .B(n6692), .Y(n1618) );
  OAI21X1 U3086 ( .A(n6502), .B(n6691), .C(n1619), .Y(n4011) );
  NAND2X1 U3087 ( .A(\Mem[53][29] ), .B(n6692), .Y(n1619) );
  OAI21X1 U3088 ( .A(n6492), .B(n6691), .C(n1620), .Y(n4012) );
  NAND2X1 U3089 ( .A(\Mem[53][30] ), .B(n6693), .Y(n1620) );
  OAI21X1 U3090 ( .A(n6487), .B(n6691), .C(n1621), .Y(n4013) );
  NAND2X1 U3091 ( .A(\Mem[53][31] ), .B(n6693), .Y(n1621) );
  NAND2X1 U3092 ( .A(n7009), .B(n7023), .Y(n1589) );
  OAI21X1 U3093 ( .A(n6607), .B(n6685), .C(n1623), .Y(n4014) );
  NAND2X1 U3094 ( .A(\Mem[54][0] ), .B(n6688), .Y(n1623) );
  OAI21X1 U3095 ( .A(n6552), .B(n6684), .C(n1624), .Y(n4015) );
  NAND2X1 U3096 ( .A(\Mem[54][1] ), .B(n6688), .Y(n1624) );
  OAI21X1 U3097 ( .A(n6497), .B(n6684), .C(n1625), .Y(n4016) );
  NAND2X1 U3098 ( .A(\Mem[54][2] ), .B(n6688), .Y(n1625) );
  OAI21X1 U3099 ( .A(n6482), .B(n6684), .C(n1626), .Y(n4017) );
  NAND2X1 U3100 ( .A(\Mem[54][3] ), .B(n6687), .Y(n1626) );
  OAI21X1 U3101 ( .A(n6477), .B(n6684), .C(n1627), .Y(n4018) );
  NAND2X1 U3102 ( .A(\Mem[54][4] ), .B(n6688), .Y(n1627) );
  OAI21X1 U3103 ( .A(n6472), .B(n6684), .C(n1628), .Y(n4019) );
  NAND2X1 U3104 ( .A(\Mem[54][5] ), .B(n6687), .Y(n1628) );
  OAI21X1 U3105 ( .A(n6467), .B(n6684), .C(n1629), .Y(n4020) );
  NAND2X1 U3106 ( .A(\Mem[54][6] ), .B(n6687), .Y(n1629) );
  OAI21X1 U3107 ( .A(n6462), .B(n6684), .C(n1630), .Y(n4021) );
  NAND2X1 U3108 ( .A(\Mem[54][7] ), .B(n6687), .Y(n1630) );
  OAI21X1 U3109 ( .A(n6457), .B(n6684), .C(n1631), .Y(n4022) );
  NAND2X1 U3110 ( .A(\Mem[54][8] ), .B(n6687), .Y(n1631) );
  OAI21X1 U3111 ( .A(n6452), .B(n6684), .C(n1632), .Y(n4023) );
  NAND2X1 U3112 ( .A(\Mem[54][9] ), .B(n6687), .Y(n1632) );
  OAI21X1 U3113 ( .A(n6602), .B(n6684), .C(n1633), .Y(n4024) );
  NAND2X1 U3114 ( .A(\Mem[54][10] ), .B(n6687), .Y(n1633) );
  OAI21X1 U3115 ( .A(n6597), .B(n6684), .C(n1634), .Y(n4025) );
  NAND2X1 U3116 ( .A(\Mem[54][11] ), .B(n6687), .Y(n1634) );
  OAI21X1 U3117 ( .A(n6592), .B(n6684), .C(n1635), .Y(n4026) );
  NAND2X1 U3118 ( .A(\Mem[54][12] ), .B(n6687), .Y(n1635) );
  OAI21X1 U3119 ( .A(n6587), .B(n6685), .C(n1636), .Y(n4027) );
  NAND2X1 U3120 ( .A(\Mem[54][13] ), .B(n6687), .Y(n1636) );
  OAI21X1 U3121 ( .A(n6582), .B(n6685), .C(n1637), .Y(n4028) );
  NAND2X1 U3122 ( .A(\Mem[54][14] ), .B(n6687), .Y(n1637) );
  OAI21X1 U3123 ( .A(n6577), .B(n6685), .C(n1638), .Y(n4029) );
  NAND2X1 U3124 ( .A(\Mem[54][15] ), .B(n6686), .Y(n1638) );
  OAI21X1 U3125 ( .A(n6572), .B(n6685), .C(n1639), .Y(n4030) );
  NAND2X1 U3126 ( .A(\Mem[54][16] ), .B(n6687), .Y(n1639) );
  OAI21X1 U3127 ( .A(n6567), .B(n6685), .C(n1640), .Y(n4031) );
  NAND2X1 U3128 ( .A(\Mem[54][17] ), .B(n6686), .Y(n1640) );
  OAI21X1 U3129 ( .A(n6562), .B(n6685), .C(n1641), .Y(n4032) );
  NAND2X1 U3130 ( .A(\Mem[54][18] ), .B(n6686), .Y(n1641) );
  OAI21X1 U3131 ( .A(n6557), .B(n6685), .C(n1642), .Y(n4033) );
  NAND2X1 U3132 ( .A(\Mem[54][19] ), .B(n6686), .Y(n1642) );
  OAI21X1 U3133 ( .A(n6547), .B(n6685), .C(n1643), .Y(n4034) );
  NAND2X1 U3134 ( .A(\Mem[54][20] ), .B(n6686), .Y(n1643) );
  OAI21X1 U3135 ( .A(n6542), .B(n6685), .C(n1644), .Y(n4035) );
  NAND2X1 U3136 ( .A(\Mem[54][21] ), .B(n6686), .Y(n1644) );
  OAI21X1 U3137 ( .A(n6537), .B(n6685), .C(n1645), .Y(n4036) );
  NAND2X1 U3138 ( .A(\Mem[54][22] ), .B(n6687), .Y(n1645) );
  OAI21X1 U3139 ( .A(n6532), .B(n6686), .C(n1646), .Y(n4037) );
  NAND2X1 U3140 ( .A(\Mem[54][23] ), .B(n6686), .Y(n1646) );
  OAI21X1 U3141 ( .A(n6527), .B(n6685), .C(n1647), .Y(n4038) );
  NAND2X1 U3142 ( .A(\Mem[54][24] ), .B(n6687), .Y(n1647) );
  OAI21X1 U3143 ( .A(n6522), .B(n6686), .C(n1648), .Y(n4039) );
  NAND2X1 U3144 ( .A(\Mem[54][25] ), .B(n6687), .Y(n1648) );
  OAI21X1 U3145 ( .A(n6517), .B(n6686), .C(n1649), .Y(n4040) );
  NAND2X1 U3146 ( .A(\Mem[54][26] ), .B(n6687), .Y(n1649) );
  OAI21X1 U3147 ( .A(n6512), .B(n6686), .C(n1650), .Y(n4041) );
  NAND2X1 U3148 ( .A(\Mem[54][27] ), .B(n6687), .Y(n1650) );
  OAI21X1 U3149 ( .A(n6507), .B(n6686), .C(n1651), .Y(n4042) );
  NAND2X1 U3150 ( .A(\Mem[54][28] ), .B(n6687), .Y(n1651) );
  OAI21X1 U3151 ( .A(n6502), .B(n6686), .C(n1652), .Y(n4043) );
  NAND2X1 U3152 ( .A(\Mem[54][29] ), .B(n6687), .Y(n1652) );
  OAI21X1 U3153 ( .A(n6492), .B(n6686), .C(n1653), .Y(n4044) );
  NAND2X1 U3154 ( .A(\Mem[54][30] ), .B(n6688), .Y(n1653) );
  OAI21X1 U3155 ( .A(n6487), .B(n6686), .C(n1654), .Y(n4045) );
  NAND2X1 U3156 ( .A(\Mem[54][31] ), .B(n6688), .Y(n1654) );
  NAND2X1 U3157 ( .A(n7009), .B(n7024), .Y(n1622) );
  OAI21X1 U3158 ( .A(n6607), .B(n6680), .C(n1656), .Y(n4046) );
  NAND2X1 U3159 ( .A(\Mem[55][0] ), .B(n6683), .Y(n1656) );
  OAI21X1 U3160 ( .A(n6552), .B(n6679), .C(n1657), .Y(n4047) );
  NAND2X1 U3161 ( .A(\Mem[55][1] ), .B(n6683), .Y(n1657) );
  OAI21X1 U3162 ( .A(n6497), .B(n6679), .C(n1658), .Y(n4048) );
  NAND2X1 U3163 ( .A(\Mem[55][2] ), .B(n6683), .Y(n1658) );
  OAI21X1 U3164 ( .A(n6482), .B(n6679), .C(n1659), .Y(n4049) );
  NAND2X1 U3165 ( .A(\Mem[55][3] ), .B(n6682), .Y(n1659) );
  OAI21X1 U3166 ( .A(n6477), .B(n6679), .C(n1660), .Y(n4050) );
  NAND2X1 U3167 ( .A(\Mem[55][4] ), .B(n6683), .Y(n1660) );
  OAI21X1 U3168 ( .A(n6472), .B(n6679), .C(n1661), .Y(n4051) );
  NAND2X1 U3169 ( .A(\Mem[55][5] ), .B(n6682), .Y(n1661) );
  OAI21X1 U3170 ( .A(n6467), .B(n6679), .C(n1662), .Y(n4052) );
  NAND2X1 U3171 ( .A(\Mem[55][6] ), .B(n6682), .Y(n1662) );
  OAI21X1 U3172 ( .A(n6462), .B(n6679), .C(n1663), .Y(n4053) );
  NAND2X1 U3173 ( .A(\Mem[55][7] ), .B(n6682), .Y(n1663) );
  OAI21X1 U3174 ( .A(n6457), .B(n6679), .C(n1664), .Y(n4054) );
  NAND2X1 U3175 ( .A(\Mem[55][8] ), .B(n6682), .Y(n1664) );
  OAI21X1 U3176 ( .A(n6452), .B(n6679), .C(n1665), .Y(n4055) );
  NAND2X1 U3177 ( .A(\Mem[55][9] ), .B(n6682), .Y(n1665) );
  OAI21X1 U3178 ( .A(n6602), .B(n6679), .C(n1666), .Y(n4056) );
  NAND2X1 U3179 ( .A(\Mem[55][10] ), .B(n6682), .Y(n1666) );
  OAI21X1 U3180 ( .A(n6597), .B(n6679), .C(n1667), .Y(n4057) );
  NAND2X1 U3181 ( .A(\Mem[55][11] ), .B(n6682), .Y(n1667) );
  OAI21X1 U3182 ( .A(n6592), .B(n6679), .C(n1668), .Y(n4058) );
  NAND2X1 U3183 ( .A(\Mem[55][12] ), .B(n6682), .Y(n1668) );
  OAI21X1 U3184 ( .A(n6587), .B(n6680), .C(n1669), .Y(n4059) );
  NAND2X1 U3185 ( .A(\Mem[55][13] ), .B(n6682), .Y(n1669) );
  OAI21X1 U3186 ( .A(n6582), .B(n6680), .C(n1670), .Y(n4060) );
  NAND2X1 U3187 ( .A(\Mem[55][14] ), .B(n6682), .Y(n1670) );
  OAI21X1 U3188 ( .A(n6577), .B(n6680), .C(n1671), .Y(n4061) );
  NAND2X1 U3189 ( .A(\Mem[55][15] ), .B(n6681), .Y(n1671) );
  OAI21X1 U3190 ( .A(n6572), .B(n6680), .C(n1672), .Y(n4062) );
  NAND2X1 U3191 ( .A(\Mem[55][16] ), .B(n6682), .Y(n1672) );
  OAI21X1 U3192 ( .A(n6567), .B(n6680), .C(n1673), .Y(n4063) );
  NAND2X1 U3193 ( .A(\Mem[55][17] ), .B(n6681), .Y(n1673) );
  OAI21X1 U3194 ( .A(n6562), .B(n6680), .C(n1674), .Y(n4064) );
  NAND2X1 U3195 ( .A(\Mem[55][18] ), .B(n6681), .Y(n1674) );
  OAI21X1 U3196 ( .A(n6557), .B(n6680), .C(n1675), .Y(n4065) );
  NAND2X1 U3197 ( .A(\Mem[55][19] ), .B(n6681), .Y(n1675) );
  OAI21X1 U3198 ( .A(n6547), .B(n6680), .C(n1676), .Y(n4066) );
  NAND2X1 U3199 ( .A(\Mem[55][20] ), .B(n6681), .Y(n1676) );
  OAI21X1 U3200 ( .A(n6542), .B(n6680), .C(n1677), .Y(n4067) );
  NAND2X1 U3201 ( .A(\Mem[55][21] ), .B(n6681), .Y(n1677) );
  OAI21X1 U3202 ( .A(n6537), .B(n6680), .C(n1678), .Y(n4068) );
  NAND2X1 U3203 ( .A(\Mem[55][22] ), .B(n6682), .Y(n1678) );
  OAI21X1 U3204 ( .A(n6532), .B(n6681), .C(n1679), .Y(n4069) );
  NAND2X1 U3205 ( .A(\Mem[55][23] ), .B(n6681), .Y(n1679) );
  OAI21X1 U3206 ( .A(n6527), .B(n6680), .C(n1680), .Y(n4070) );
  NAND2X1 U3207 ( .A(\Mem[55][24] ), .B(n6682), .Y(n1680) );
  OAI21X1 U3208 ( .A(n6522), .B(n6681), .C(n1681), .Y(n4071) );
  NAND2X1 U3209 ( .A(\Mem[55][25] ), .B(n6682), .Y(n1681) );
  OAI21X1 U3210 ( .A(n6517), .B(n6681), .C(n1682), .Y(n4072) );
  NAND2X1 U3211 ( .A(\Mem[55][26] ), .B(n6682), .Y(n1682) );
  OAI21X1 U3212 ( .A(n6512), .B(n6681), .C(n1683), .Y(n4073) );
  NAND2X1 U3213 ( .A(\Mem[55][27] ), .B(n6682), .Y(n1683) );
  OAI21X1 U3214 ( .A(n6507), .B(n6681), .C(n1684), .Y(n4074) );
  NAND2X1 U3215 ( .A(\Mem[55][28] ), .B(n6682), .Y(n1684) );
  OAI21X1 U3216 ( .A(n6502), .B(n6681), .C(n1685), .Y(n4075) );
  NAND2X1 U3217 ( .A(\Mem[55][29] ), .B(n6682), .Y(n1685) );
  OAI21X1 U3218 ( .A(n6492), .B(n6681), .C(n1686), .Y(n4076) );
  NAND2X1 U3219 ( .A(\Mem[55][30] ), .B(n6683), .Y(n1686) );
  OAI21X1 U3220 ( .A(n6487), .B(n6681), .C(n1687), .Y(n4077) );
  NAND2X1 U3221 ( .A(\Mem[55][31] ), .B(n6683), .Y(n1687) );
  NAND2X1 U3222 ( .A(n7009), .B(n7021), .Y(n1655) );
  NAND3X1 U3224 ( .A(ADDR_WR[4]), .B(n7015), .C(n80), .Y(n1688) );
  OAI21X1 U3225 ( .A(n6607), .B(n6675), .C(n1690), .Y(n4078) );
  NAND2X1 U3226 ( .A(\Mem[56][0] ), .B(n6678), .Y(n1690) );
  OAI21X1 U3227 ( .A(n6552), .B(n6674), .C(n1691), .Y(n4079) );
  NAND2X1 U3228 ( .A(\Mem[56][1] ), .B(n6678), .Y(n1691) );
  OAI21X1 U3229 ( .A(n6497), .B(n6674), .C(n1692), .Y(n4080) );
  NAND2X1 U3230 ( .A(\Mem[56][2] ), .B(n6678), .Y(n1692) );
  OAI21X1 U3231 ( .A(n6482), .B(n6674), .C(n1693), .Y(n4081) );
  NAND2X1 U3232 ( .A(\Mem[56][3] ), .B(n6677), .Y(n1693) );
  OAI21X1 U3233 ( .A(n6477), .B(n6674), .C(n1694), .Y(n4082) );
  NAND2X1 U3234 ( .A(\Mem[56][4] ), .B(n6678), .Y(n1694) );
  OAI21X1 U3235 ( .A(n6472), .B(n6674), .C(n1695), .Y(n4083) );
  NAND2X1 U3236 ( .A(\Mem[56][5] ), .B(n6677), .Y(n1695) );
  OAI21X1 U3237 ( .A(n6467), .B(n6674), .C(n1696), .Y(n4084) );
  NAND2X1 U3238 ( .A(\Mem[56][6] ), .B(n6677), .Y(n1696) );
  OAI21X1 U3239 ( .A(n6462), .B(n6674), .C(n1697), .Y(n4085) );
  NAND2X1 U3240 ( .A(\Mem[56][7] ), .B(n6677), .Y(n1697) );
  OAI21X1 U3241 ( .A(n6457), .B(n6674), .C(n1698), .Y(n4086) );
  NAND2X1 U3242 ( .A(\Mem[56][8] ), .B(n6677), .Y(n1698) );
  OAI21X1 U3243 ( .A(n6452), .B(n6674), .C(n1699), .Y(n4087) );
  NAND2X1 U3244 ( .A(\Mem[56][9] ), .B(n6677), .Y(n1699) );
  OAI21X1 U3245 ( .A(n6602), .B(n6674), .C(n1700), .Y(n4088) );
  NAND2X1 U3246 ( .A(\Mem[56][10] ), .B(n6677), .Y(n1700) );
  OAI21X1 U3247 ( .A(n6597), .B(n6674), .C(n1701), .Y(n4089) );
  NAND2X1 U3248 ( .A(\Mem[56][11] ), .B(n6677), .Y(n1701) );
  OAI21X1 U3249 ( .A(n6592), .B(n6674), .C(n1702), .Y(n4090) );
  NAND2X1 U3250 ( .A(\Mem[56][12] ), .B(n6677), .Y(n1702) );
  OAI21X1 U3251 ( .A(n6587), .B(n6675), .C(n1703), .Y(n4091) );
  NAND2X1 U3252 ( .A(\Mem[56][13] ), .B(n6677), .Y(n1703) );
  OAI21X1 U3253 ( .A(n6582), .B(n6675), .C(n1704), .Y(n4092) );
  NAND2X1 U3254 ( .A(\Mem[56][14] ), .B(n6677), .Y(n1704) );
  OAI21X1 U3255 ( .A(n6577), .B(n6675), .C(n1705), .Y(n4093) );
  NAND2X1 U3256 ( .A(\Mem[56][15] ), .B(n6676), .Y(n1705) );
  OAI21X1 U3257 ( .A(n6572), .B(n6675), .C(n1706), .Y(n4094) );
  NAND2X1 U3258 ( .A(\Mem[56][16] ), .B(n6677), .Y(n1706) );
  OAI21X1 U3259 ( .A(n6567), .B(n6675), .C(n1707), .Y(n4095) );
  NAND2X1 U3260 ( .A(\Mem[56][17] ), .B(n6676), .Y(n1707) );
  OAI21X1 U3261 ( .A(n6562), .B(n6675), .C(n1708), .Y(n4096) );
  NAND2X1 U3262 ( .A(\Mem[56][18] ), .B(n6676), .Y(n1708) );
  OAI21X1 U3263 ( .A(n6557), .B(n6675), .C(n1709), .Y(n4097) );
  NAND2X1 U3264 ( .A(\Mem[56][19] ), .B(n6676), .Y(n1709) );
  OAI21X1 U3265 ( .A(n6547), .B(n6675), .C(n1710), .Y(n4098) );
  NAND2X1 U3266 ( .A(\Mem[56][20] ), .B(n6676), .Y(n1710) );
  OAI21X1 U3267 ( .A(n6542), .B(n6675), .C(n1711), .Y(n4099) );
  NAND2X1 U3268 ( .A(\Mem[56][21] ), .B(n6676), .Y(n1711) );
  OAI21X1 U3269 ( .A(n6537), .B(n6675), .C(n1712), .Y(n4100) );
  NAND2X1 U3270 ( .A(\Mem[56][22] ), .B(n6677), .Y(n1712) );
  OAI21X1 U3271 ( .A(n6532), .B(n6676), .C(n1713), .Y(n4101) );
  NAND2X1 U3272 ( .A(\Mem[56][23] ), .B(n6676), .Y(n1713) );
  OAI21X1 U3273 ( .A(n6527), .B(n6675), .C(n1714), .Y(n4102) );
  NAND2X1 U3274 ( .A(\Mem[56][24] ), .B(n6677), .Y(n1714) );
  OAI21X1 U3275 ( .A(n6522), .B(n6676), .C(n1715), .Y(n4103) );
  NAND2X1 U3276 ( .A(\Mem[56][25] ), .B(n6677), .Y(n1715) );
  OAI21X1 U3277 ( .A(n6517), .B(n6676), .C(n1716), .Y(n4104) );
  NAND2X1 U3278 ( .A(\Mem[56][26] ), .B(n6677), .Y(n1716) );
  OAI21X1 U3279 ( .A(n6512), .B(n6676), .C(n1717), .Y(n4105) );
  NAND2X1 U3280 ( .A(\Mem[56][27] ), .B(n6677), .Y(n1717) );
  OAI21X1 U3281 ( .A(n6507), .B(n6676), .C(n1718), .Y(n4106) );
  NAND2X1 U3282 ( .A(\Mem[56][28] ), .B(n6677), .Y(n1718) );
  OAI21X1 U3283 ( .A(n6502), .B(n6676), .C(n1719), .Y(n4107) );
  NAND2X1 U3284 ( .A(\Mem[56][29] ), .B(n6677), .Y(n1719) );
  OAI21X1 U3285 ( .A(n6492), .B(n6676), .C(n1720), .Y(n4108) );
  NAND2X1 U3286 ( .A(\Mem[56][30] ), .B(n6678), .Y(n1720) );
  OAI21X1 U3287 ( .A(n6487), .B(n6676), .C(n1721), .Y(n4109) );
  NAND2X1 U3288 ( .A(\Mem[56][31] ), .B(n6678), .Y(n1721) );
  NAND2X1 U3289 ( .A(n7008), .B(n7016), .Y(n1689) );
  OAI21X1 U3290 ( .A(n6608), .B(n6670), .C(n1724), .Y(n4110) );
  NAND2X1 U3291 ( .A(\Mem[57][0] ), .B(n6673), .Y(n1724) );
  OAI21X1 U3292 ( .A(n6553), .B(n6669), .C(n1725), .Y(n4111) );
  NAND2X1 U3293 ( .A(\Mem[57][1] ), .B(n6673), .Y(n1725) );
  OAI21X1 U3294 ( .A(n6498), .B(n6669), .C(n1726), .Y(n4112) );
  NAND2X1 U3295 ( .A(\Mem[57][2] ), .B(n6673), .Y(n1726) );
  OAI21X1 U3296 ( .A(n6483), .B(n6669), .C(n1727), .Y(n4113) );
  NAND2X1 U3297 ( .A(\Mem[57][3] ), .B(n6672), .Y(n1727) );
  OAI21X1 U3298 ( .A(n6478), .B(n6669), .C(n1728), .Y(n4114) );
  NAND2X1 U3299 ( .A(\Mem[57][4] ), .B(n6673), .Y(n1728) );
  OAI21X1 U3300 ( .A(n6473), .B(n6669), .C(n1729), .Y(n4115) );
  NAND2X1 U3301 ( .A(\Mem[57][5] ), .B(n6672), .Y(n1729) );
  OAI21X1 U3302 ( .A(n6468), .B(n6669), .C(n1730), .Y(n4116) );
  NAND2X1 U3303 ( .A(\Mem[57][6] ), .B(n6672), .Y(n1730) );
  OAI21X1 U3304 ( .A(n6463), .B(n6669), .C(n1731), .Y(n4117) );
  NAND2X1 U3305 ( .A(\Mem[57][7] ), .B(n6672), .Y(n1731) );
  OAI21X1 U3306 ( .A(n6458), .B(n6669), .C(n1732), .Y(n4118) );
  NAND2X1 U3307 ( .A(\Mem[57][8] ), .B(n6672), .Y(n1732) );
  OAI21X1 U3308 ( .A(n6453), .B(n6669), .C(n1733), .Y(n4119) );
  NAND2X1 U3309 ( .A(\Mem[57][9] ), .B(n6672), .Y(n1733) );
  OAI21X1 U3310 ( .A(n6603), .B(n6669), .C(n1734), .Y(n4120) );
  NAND2X1 U3311 ( .A(\Mem[57][10] ), .B(n6672), .Y(n1734) );
  OAI21X1 U3312 ( .A(n6598), .B(n6669), .C(n1735), .Y(n4121) );
  NAND2X1 U3313 ( .A(\Mem[57][11] ), .B(n6672), .Y(n1735) );
  OAI21X1 U3314 ( .A(n6593), .B(n6669), .C(n1736), .Y(n4122) );
  NAND2X1 U3315 ( .A(\Mem[57][12] ), .B(n6672), .Y(n1736) );
  OAI21X1 U3316 ( .A(n6588), .B(n6670), .C(n1737), .Y(n4123) );
  NAND2X1 U3317 ( .A(\Mem[57][13] ), .B(n6672), .Y(n1737) );
  OAI21X1 U3318 ( .A(n6583), .B(n6670), .C(n1738), .Y(n4124) );
  NAND2X1 U3319 ( .A(\Mem[57][14] ), .B(n6672), .Y(n1738) );
  OAI21X1 U3320 ( .A(n6578), .B(n6670), .C(n1739), .Y(n4125) );
  NAND2X1 U3321 ( .A(\Mem[57][15] ), .B(n6671), .Y(n1739) );
  OAI21X1 U3322 ( .A(n6573), .B(n6670), .C(n1740), .Y(n4126) );
  NAND2X1 U3323 ( .A(\Mem[57][16] ), .B(n6672), .Y(n1740) );
  OAI21X1 U3324 ( .A(n6568), .B(n6670), .C(n1741), .Y(n4127) );
  NAND2X1 U3325 ( .A(\Mem[57][17] ), .B(n6671), .Y(n1741) );
  OAI21X1 U3326 ( .A(n6563), .B(n6670), .C(n1742), .Y(n4128) );
  NAND2X1 U3327 ( .A(\Mem[57][18] ), .B(n6671), .Y(n1742) );
  OAI21X1 U3328 ( .A(n6557), .B(n6670), .C(n1743), .Y(n4129) );
  NAND2X1 U3329 ( .A(\Mem[57][19] ), .B(n6671), .Y(n1743) );
  OAI21X1 U3330 ( .A(n6547), .B(n6670), .C(n1744), .Y(n4130) );
  NAND2X1 U3331 ( .A(\Mem[57][20] ), .B(n6671), .Y(n1744) );
  OAI21X1 U3332 ( .A(n6542), .B(n6670), .C(n1745), .Y(n4131) );
  NAND2X1 U3333 ( .A(\Mem[57][21] ), .B(n6671), .Y(n1745) );
  OAI21X1 U3334 ( .A(n6537), .B(n6670), .C(n1746), .Y(n4132) );
  NAND2X1 U3335 ( .A(\Mem[57][22] ), .B(n6672), .Y(n1746) );
  OAI21X1 U3336 ( .A(n6532), .B(n6671), .C(n1747), .Y(n4133) );
  NAND2X1 U3337 ( .A(\Mem[57][23] ), .B(n6671), .Y(n1747) );
  OAI21X1 U3338 ( .A(n6527), .B(n6670), .C(n1748), .Y(n4134) );
  NAND2X1 U3339 ( .A(\Mem[57][24] ), .B(n6672), .Y(n1748) );
  OAI21X1 U3340 ( .A(n6522), .B(n6671), .C(n1749), .Y(n4135) );
  NAND2X1 U3341 ( .A(\Mem[57][25] ), .B(n6672), .Y(n1749) );
  OAI21X1 U3342 ( .A(n6517), .B(n6671), .C(n1750), .Y(n4136) );
  NAND2X1 U3343 ( .A(\Mem[57][26] ), .B(n6672), .Y(n1750) );
  OAI21X1 U3344 ( .A(n6512), .B(n6671), .C(n1751), .Y(n4137) );
  NAND2X1 U3345 ( .A(\Mem[57][27] ), .B(n6672), .Y(n1751) );
  OAI21X1 U3346 ( .A(n6507), .B(n6671), .C(n1752), .Y(n4138) );
  NAND2X1 U3347 ( .A(\Mem[57][28] ), .B(n6672), .Y(n1752) );
  OAI21X1 U3348 ( .A(n6502), .B(n6671), .C(n1753), .Y(n4139) );
  NAND2X1 U3349 ( .A(\Mem[57][29] ), .B(n6672), .Y(n1753) );
  OAI21X1 U3350 ( .A(n6492), .B(n6671), .C(n1754), .Y(n4140) );
  NAND2X1 U3351 ( .A(\Mem[57][30] ), .B(n6673), .Y(n1754) );
  OAI21X1 U3352 ( .A(n6487), .B(n6671), .C(n1755), .Y(n4141) );
  NAND2X1 U3353 ( .A(\Mem[57][31] ), .B(n6673), .Y(n1755) );
  NAND2X1 U3354 ( .A(n7008), .B(n7017), .Y(n1723) );
  OAI21X1 U3355 ( .A(n6608), .B(n6665), .C(n1757), .Y(n4142) );
  NAND2X1 U3356 ( .A(\Mem[58][0] ), .B(n6668), .Y(n1757) );
  OAI21X1 U3357 ( .A(n6553), .B(n6664), .C(n1758), .Y(n4143) );
  NAND2X1 U3358 ( .A(\Mem[58][1] ), .B(n6668), .Y(n1758) );
  OAI21X1 U3359 ( .A(n6498), .B(n6664), .C(n1759), .Y(n4144) );
  NAND2X1 U3360 ( .A(\Mem[58][2] ), .B(n6668), .Y(n1759) );
  OAI21X1 U3361 ( .A(n6483), .B(n6664), .C(n1760), .Y(n4145) );
  NAND2X1 U3362 ( .A(\Mem[58][3] ), .B(n6667), .Y(n1760) );
  OAI21X1 U3363 ( .A(n6478), .B(n6664), .C(n1761), .Y(n4146) );
  NAND2X1 U3364 ( .A(\Mem[58][4] ), .B(n6668), .Y(n1761) );
  OAI21X1 U3365 ( .A(n6473), .B(n6664), .C(n1762), .Y(n4147) );
  NAND2X1 U3366 ( .A(\Mem[58][5] ), .B(n6667), .Y(n1762) );
  OAI21X1 U3367 ( .A(n6468), .B(n6664), .C(n1763), .Y(n4148) );
  NAND2X1 U3368 ( .A(\Mem[58][6] ), .B(n6667), .Y(n1763) );
  OAI21X1 U3369 ( .A(n6463), .B(n6664), .C(n1764), .Y(n4149) );
  NAND2X1 U3370 ( .A(\Mem[58][7] ), .B(n6667), .Y(n1764) );
  OAI21X1 U3371 ( .A(n6458), .B(n6664), .C(n1765), .Y(n4150) );
  NAND2X1 U3372 ( .A(\Mem[58][8] ), .B(n6667), .Y(n1765) );
  OAI21X1 U3373 ( .A(n6453), .B(n6664), .C(n1766), .Y(n4151) );
  NAND2X1 U3374 ( .A(\Mem[58][9] ), .B(n6667), .Y(n1766) );
  OAI21X1 U3375 ( .A(n6603), .B(n6664), .C(n1767), .Y(n4152) );
  NAND2X1 U3376 ( .A(\Mem[58][10] ), .B(n6667), .Y(n1767) );
  OAI21X1 U3377 ( .A(n6598), .B(n6664), .C(n1768), .Y(n4153) );
  NAND2X1 U3378 ( .A(\Mem[58][11] ), .B(n6667), .Y(n1768) );
  OAI21X1 U3379 ( .A(n6593), .B(n6664), .C(n1769), .Y(n4154) );
  NAND2X1 U3380 ( .A(\Mem[58][12] ), .B(n6667), .Y(n1769) );
  OAI21X1 U3381 ( .A(n6588), .B(n6665), .C(n1770), .Y(n4155) );
  NAND2X1 U3382 ( .A(\Mem[58][13] ), .B(n6667), .Y(n1770) );
  OAI21X1 U3383 ( .A(n6583), .B(n6665), .C(n1771), .Y(n4156) );
  NAND2X1 U3384 ( .A(\Mem[58][14] ), .B(n6667), .Y(n1771) );
  OAI21X1 U3385 ( .A(n6578), .B(n6665), .C(n1772), .Y(n4157) );
  NAND2X1 U3386 ( .A(\Mem[58][15] ), .B(n6666), .Y(n1772) );
  OAI21X1 U3387 ( .A(n6573), .B(n6665), .C(n1773), .Y(n4158) );
  NAND2X1 U3388 ( .A(\Mem[58][16] ), .B(n6667), .Y(n1773) );
  OAI21X1 U3389 ( .A(n6568), .B(n6665), .C(n1774), .Y(n4159) );
  NAND2X1 U3390 ( .A(\Mem[58][17] ), .B(n6666), .Y(n1774) );
  OAI21X1 U3391 ( .A(n6563), .B(n6665), .C(n1775), .Y(n4160) );
  NAND2X1 U3392 ( .A(\Mem[58][18] ), .B(n6666), .Y(n1775) );
  OAI21X1 U3393 ( .A(n6558), .B(n6665), .C(n1776), .Y(n4161) );
  NAND2X1 U3394 ( .A(\Mem[58][19] ), .B(n6666), .Y(n1776) );
  OAI21X1 U3395 ( .A(n6548), .B(n6665), .C(n1777), .Y(n4162) );
  NAND2X1 U3396 ( .A(\Mem[58][20] ), .B(n6666), .Y(n1777) );
  OAI21X1 U3397 ( .A(n6543), .B(n6665), .C(n1778), .Y(n4163) );
  NAND2X1 U3398 ( .A(\Mem[58][21] ), .B(n6666), .Y(n1778) );
  OAI21X1 U3399 ( .A(n6538), .B(n6665), .C(n1779), .Y(n4164) );
  NAND2X1 U3400 ( .A(\Mem[58][22] ), .B(n6667), .Y(n1779) );
  OAI21X1 U3401 ( .A(n6533), .B(n6666), .C(n1780), .Y(n4165) );
  NAND2X1 U3402 ( .A(\Mem[58][23] ), .B(n6666), .Y(n1780) );
  OAI21X1 U3403 ( .A(n6528), .B(n6665), .C(n1781), .Y(n4166) );
  NAND2X1 U3404 ( .A(\Mem[58][24] ), .B(n6667), .Y(n1781) );
  OAI21X1 U3405 ( .A(n6523), .B(n6666), .C(n1782), .Y(n4167) );
  NAND2X1 U3406 ( .A(\Mem[58][25] ), .B(n6667), .Y(n1782) );
  OAI21X1 U3407 ( .A(n6518), .B(n6666), .C(n1783), .Y(n4168) );
  NAND2X1 U3408 ( .A(\Mem[58][26] ), .B(n6667), .Y(n1783) );
  OAI21X1 U3409 ( .A(n6513), .B(n6666), .C(n1784), .Y(n4169) );
  NAND2X1 U3410 ( .A(\Mem[58][27] ), .B(n6667), .Y(n1784) );
  OAI21X1 U3411 ( .A(n6508), .B(n6666), .C(n1785), .Y(n4170) );
  NAND2X1 U3412 ( .A(\Mem[58][28] ), .B(n6667), .Y(n1785) );
  OAI21X1 U3413 ( .A(n6503), .B(n6666), .C(n1786), .Y(n4171) );
  NAND2X1 U3414 ( .A(\Mem[58][29] ), .B(n6667), .Y(n1786) );
  OAI21X1 U3415 ( .A(n6493), .B(n6666), .C(n1787), .Y(n4172) );
  NAND2X1 U3416 ( .A(\Mem[58][30] ), .B(n6668), .Y(n1787) );
  OAI21X1 U3417 ( .A(n6488), .B(n6666), .C(n1788), .Y(n4173) );
  NAND2X1 U3418 ( .A(\Mem[58][31] ), .B(n6668), .Y(n1788) );
  NAND2X1 U3419 ( .A(n7008), .B(n7018), .Y(n1756) );
  OAI21X1 U3420 ( .A(n6608), .B(n6660), .C(n1790), .Y(n4174) );
  NAND2X1 U3421 ( .A(\Mem[59][0] ), .B(n6663), .Y(n1790) );
  OAI21X1 U3422 ( .A(n6553), .B(n6659), .C(n1791), .Y(n4175) );
  NAND2X1 U3423 ( .A(\Mem[59][1] ), .B(n6663), .Y(n1791) );
  OAI21X1 U3424 ( .A(n6498), .B(n6659), .C(n1792), .Y(n4176) );
  NAND2X1 U3425 ( .A(\Mem[59][2] ), .B(n6663), .Y(n1792) );
  OAI21X1 U3426 ( .A(n6483), .B(n6659), .C(n1793), .Y(n4177) );
  NAND2X1 U3427 ( .A(\Mem[59][3] ), .B(n6662), .Y(n1793) );
  OAI21X1 U3428 ( .A(n6478), .B(n6659), .C(n1794), .Y(n4178) );
  NAND2X1 U3429 ( .A(\Mem[59][4] ), .B(n6663), .Y(n1794) );
  OAI21X1 U3430 ( .A(n6473), .B(n6659), .C(n1795), .Y(n4179) );
  NAND2X1 U3431 ( .A(\Mem[59][5] ), .B(n6662), .Y(n1795) );
  OAI21X1 U3432 ( .A(n6468), .B(n6659), .C(n1796), .Y(n4180) );
  NAND2X1 U3433 ( .A(\Mem[59][6] ), .B(n6662), .Y(n1796) );
  OAI21X1 U3434 ( .A(n6463), .B(n6659), .C(n1797), .Y(n4181) );
  NAND2X1 U3435 ( .A(\Mem[59][7] ), .B(n6662), .Y(n1797) );
  OAI21X1 U3436 ( .A(n6458), .B(n6659), .C(n1798), .Y(n4182) );
  NAND2X1 U3437 ( .A(\Mem[59][8] ), .B(n6662), .Y(n1798) );
  OAI21X1 U3438 ( .A(n6453), .B(n6659), .C(n1799), .Y(n4183) );
  NAND2X1 U3439 ( .A(\Mem[59][9] ), .B(n6662), .Y(n1799) );
  OAI21X1 U3440 ( .A(n6603), .B(n6659), .C(n1800), .Y(n4184) );
  NAND2X1 U3441 ( .A(\Mem[59][10] ), .B(n6662), .Y(n1800) );
  OAI21X1 U3442 ( .A(n6598), .B(n6659), .C(n1801), .Y(n4185) );
  NAND2X1 U3443 ( .A(\Mem[59][11] ), .B(n6662), .Y(n1801) );
  OAI21X1 U3444 ( .A(n6593), .B(n6659), .C(n1802), .Y(n4186) );
  NAND2X1 U3445 ( .A(\Mem[59][12] ), .B(n6662), .Y(n1802) );
  OAI21X1 U3446 ( .A(n6588), .B(n6660), .C(n1803), .Y(n4187) );
  NAND2X1 U3447 ( .A(\Mem[59][13] ), .B(n6662), .Y(n1803) );
  OAI21X1 U3448 ( .A(n6583), .B(n6660), .C(n1804), .Y(n4188) );
  NAND2X1 U3449 ( .A(\Mem[59][14] ), .B(n6662), .Y(n1804) );
  OAI21X1 U3450 ( .A(n6578), .B(n6660), .C(n1805), .Y(n4189) );
  NAND2X1 U3451 ( .A(\Mem[59][15] ), .B(n6661), .Y(n1805) );
  OAI21X1 U3452 ( .A(n6573), .B(n6660), .C(n1806), .Y(n4190) );
  NAND2X1 U3453 ( .A(\Mem[59][16] ), .B(n6662), .Y(n1806) );
  OAI21X1 U3454 ( .A(n6568), .B(n6660), .C(n1807), .Y(n4191) );
  NAND2X1 U3455 ( .A(\Mem[59][17] ), .B(n6661), .Y(n1807) );
  OAI21X1 U3456 ( .A(n6563), .B(n6660), .C(n1808), .Y(n4192) );
  NAND2X1 U3457 ( .A(\Mem[59][18] ), .B(n6661), .Y(n1808) );
  OAI21X1 U3458 ( .A(n6558), .B(n6660), .C(n1809), .Y(n4193) );
  NAND2X1 U3459 ( .A(\Mem[59][19] ), .B(n6661), .Y(n1809) );
  OAI21X1 U3460 ( .A(n6548), .B(n6660), .C(n1810), .Y(n4194) );
  NAND2X1 U3461 ( .A(\Mem[59][20] ), .B(n6661), .Y(n1810) );
  OAI21X1 U3462 ( .A(n6543), .B(n6660), .C(n1811), .Y(n4195) );
  NAND2X1 U3463 ( .A(\Mem[59][21] ), .B(n6661), .Y(n1811) );
  OAI21X1 U3464 ( .A(n6538), .B(n6660), .C(n1812), .Y(n4196) );
  NAND2X1 U3465 ( .A(\Mem[59][22] ), .B(n6662), .Y(n1812) );
  OAI21X1 U3466 ( .A(n6533), .B(n6661), .C(n1813), .Y(n4197) );
  NAND2X1 U3467 ( .A(\Mem[59][23] ), .B(n6661), .Y(n1813) );
  OAI21X1 U3468 ( .A(n6528), .B(n6660), .C(n1814), .Y(n4198) );
  NAND2X1 U3469 ( .A(\Mem[59][24] ), .B(n6662), .Y(n1814) );
  OAI21X1 U3470 ( .A(n6523), .B(n6661), .C(n1815), .Y(n4199) );
  NAND2X1 U3471 ( .A(\Mem[59][25] ), .B(n6662), .Y(n1815) );
  OAI21X1 U3472 ( .A(n6518), .B(n6661), .C(n1816), .Y(n4200) );
  NAND2X1 U3473 ( .A(\Mem[59][26] ), .B(n6662), .Y(n1816) );
  OAI21X1 U3474 ( .A(n6513), .B(n6661), .C(n1817), .Y(n4201) );
  NAND2X1 U3475 ( .A(\Mem[59][27] ), .B(n6662), .Y(n1817) );
  OAI21X1 U3476 ( .A(n6508), .B(n6661), .C(n1818), .Y(n4202) );
  NAND2X1 U3477 ( .A(\Mem[59][28] ), .B(n6662), .Y(n1818) );
  OAI21X1 U3478 ( .A(n6503), .B(n6661), .C(n1819), .Y(n4203) );
  NAND2X1 U3479 ( .A(\Mem[59][29] ), .B(n6662), .Y(n1819) );
  OAI21X1 U3480 ( .A(n6493), .B(n6661), .C(n1820), .Y(n4204) );
  NAND2X1 U3481 ( .A(\Mem[59][30] ), .B(n6663), .Y(n1820) );
  OAI21X1 U3482 ( .A(n6488), .B(n6661), .C(n1821), .Y(n4205) );
  NAND2X1 U3483 ( .A(\Mem[59][31] ), .B(n6663), .Y(n1821) );
  NAND2X1 U3484 ( .A(n7008), .B(n7019), .Y(n1789) );
  OAI21X1 U3485 ( .A(n6608), .B(n6655), .C(n1823), .Y(n4206) );
  NAND2X1 U3486 ( .A(\Mem[60][0] ), .B(n6658), .Y(n1823) );
  OAI21X1 U3487 ( .A(n6553), .B(n6654), .C(n1824), .Y(n4207) );
  NAND2X1 U3488 ( .A(\Mem[60][1] ), .B(n6658), .Y(n1824) );
  OAI21X1 U3489 ( .A(n6498), .B(n6654), .C(n1825), .Y(n4208) );
  NAND2X1 U3490 ( .A(\Mem[60][2] ), .B(n6658), .Y(n1825) );
  OAI21X1 U3491 ( .A(n6483), .B(n6654), .C(n1826), .Y(n4209) );
  NAND2X1 U3492 ( .A(\Mem[60][3] ), .B(n6657), .Y(n1826) );
  OAI21X1 U3493 ( .A(n6478), .B(n6654), .C(n1827), .Y(n4210) );
  NAND2X1 U3494 ( .A(\Mem[60][4] ), .B(n6658), .Y(n1827) );
  OAI21X1 U3495 ( .A(n6473), .B(n6654), .C(n1828), .Y(n4211) );
  NAND2X1 U3496 ( .A(\Mem[60][5] ), .B(n6657), .Y(n1828) );
  OAI21X1 U3497 ( .A(n6468), .B(n6654), .C(n1829), .Y(n4212) );
  NAND2X1 U3498 ( .A(\Mem[60][6] ), .B(n6657), .Y(n1829) );
  OAI21X1 U3499 ( .A(n6463), .B(n6654), .C(n1830), .Y(n4213) );
  NAND2X1 U3500 ( .A(\Mem[60][7] ), .B(n6657), .Y(n1830) );
  OAI21X1 U3501 ( .A(n6458), .B(n6654), .C(n1831), .Y(n4214) );
  NAND2X1 U3502 ( .A(\Mem[60][8] ), .B(n6657), .Y(n1831) );
  OAI21X1 U3503 ( .A(n6453), .B(n6654), .C(n1832), .Y(n4215) );
  NAND2X1 U3504 ( .A(\Mem[60][9] ), .B(n6657), .Y(n1832) );
  OAI21X1 U3505 ( .A(n6603), .B(n6654), .C(n1833), .Y(n4216) );
  NAND2X1 U3506 ( .A(\Mem[60][10] ), .B(n6657), .Y(n1833) );
  OAI21X1 U3507 ( .A(n6598), .B(n6654), .C(n1834), .Y(n4217) );
  NAND2X1 U3508 ( .A(\Mem[60][11] ), .B(n6657), .Y(n1834) );
  OAI21X1 U3509 ( .A(n6593), .B(n6654), .C(n1835), .Y(n4218) );
  NAND2X1 U3510 ( .A(\Mem[60][12] ), .B(n6657), .Y(n1835) );
  OAI21X1 U3511 ( .A(n6588), .B(n6655), .C(n1836), .Y(n4219) );
  NAND2X1 U3512 ( .A(\Mem[60][13] ), .B(n6657), .Y(n1836) );
  OAI21X1 U3513 ( .A(n6583), .B(n6655), .C(n1837), .Y(n4220) );
  NAND2X1 U3514 ( .A(\Mem[60][14] ), .B(n6657), .Y(n1837) );
  OAI21X1 U3515 ( .A(n6578), .B(n6655), .C(n1838), .Y(n4221) );
  NAND2X1 U3516 ( .A(\Mem[60][15] ), .B(n6656), .Y(n1838) );
  OAI21X1 U3517 ( .A(n6573), .B(n6655), .C(n1839), .Y(n4222) );
  NAND2X1 U3518 ( .A(\Mem[60][16] ), .B(n6657), .Y(n1839) );
  OAI21X1 U3519 ( .A(n6568), .B(n6655), .C(n1840), .Y(n4223) );
  NAND2X1 U3520 ( .A(\Mem[60][17] ), .B(n6656), .Y(n1840) );
  OAI21X1 U3521 ( .A(n6563), .B(n6655), .C(n1841), .Y(n4224) );
  NAND2X1 U3522 ( .A(\Mem[60][18] ), .B(n6656), .Y(n1841) );
  OAI21X1 U3523 ( .A(n6558), .B(n6655), .C(n1842), .Y(n4225) );
  NAND2X1 U3524 ( .A(\Mem[60][19] ), .B(n6656), .Y(n1842) );
  OAI21X1 U3525 ( .A(n6548), .B(n6655), .C(n1843), .Y(n4226) );
  NAND2X1 U3526 ( .A(\Mem[60][20] ), .B(n6656), .Y(n1843) );
  OAI21X1 U3527 ( .A(n6543), .B(n6655), .C(n1844), .Y(n4227) );
  NAND2X1 U3528 ( .A(\Mem[60][21] ), .B(n6656), .Y(n1844) );
  OAI21X1 U3529 ( .A(n6538), .B(n6655), .C(n1845), .Y(n4228) );
  NAND2X1 U3530 ( .A(\Mem[60][22] ), .B(n6657), .Y(n1845) );
  OAI21X1 U3531 ( .A(n6533), .B(n6656), .C(n1846), .Y(n4229) );
  NAND2X1 U3532 ( .A(\Mem[60][23] ), .B(n6656), .Y(n1846) );
  OAI21X1 U3533 ( .A(n6528), .B(n6655), .C(n1847), .Y(n4230) );
  NAND2X1 U3534 ( .A(\Mem[60][24] ), .B(n6657), .Y(n1847) );
  OAI21X1 U3535 ( .A(n6523), .B(n6656), .C(n1848), .Y(n4231) );
  NAND2X1 U3536 ( .A(\Mem[60][25] ), .B(n6657), .Y(n1848) );
  OAI21X1 U3537 ( .A(n6518), .B(n6656), .C(n1849), .Y(n4232) );
  NAND2X1 U3538 ( .A(\Mem[60][26] ), .B(n6657), .Y(n1849) );
  OAI21X1 U3539 ( .A(n6513), .B(n6656), .C(n1850), .Y(n4233) );
  NAND2X1 U3540 ( .A(\Mem[60][27] ), .B(n6657), .Y(n1850) );
  OAI21X1 U3541 ( .A(n6508), .B(n6656), .C(n1851), .Y(n4234) );
  NAND2X1 U3542 ( .A(\Mem[60][28] ), .B(n6657), .Y(n1851) );
  OAI21X1 U3543 ( .A(n6503), .B(n6656), .C(n1852), .Y(n4235) );
  NAND2X1 U3544 ( .A(\Mem[60][29] ), .B(n6657), .Y(n1852) );
  OAI21X1 U3545 ( .A(n6493), .B(n6656), .C(n1853), .Y(n4236) );
  NAND2X1 U3546 ( .A(\Mem[60][30] ), .B(n6658), .Y(n1853) );
  OAI21X1 U3547 ( .A(n6488), .B(n6656), .C(n1854), .Y(n4237) );
  NAND2X1 U3548 ( .A(\Mem[60][31] ), .B(n6658), .Y(n1854) );
  NAND2X1 U3549 ( .A(n7008), .B(n7022), .Y(n1822) );
  OAI21X1 U3550 ( .A(n6608), .B(n6650), .C(n1856), .Y(n4238) );
  NAND2X1 U3551 ( .A(\Mem[61][0] ), .B(n6653), .Y(n1856) );
  OAI21X1 U3552 ( .A(n6553), .B(n6649), .C(n1857), .Y(n4239) );
  NAND2X1 U3553 ( .A(\Mem[61][1] ), .B(n6653), .Y(n1857) );
  OAI21X1 U3554 ( .A(n6498), .B(n6649), .C(n1858), .Y(n4240) );
  NAND2X1 U3555 ( .A(\Mem[61][2] ), .B(n6653), .Y(n1858) );
  OAI21X1 U3556 ( .A(n6483), .B(n6649), .C(n1859), .Y(n4241) );
  NAND2X1 U3557 ( .A(\Mem[61][3] ), .B(n6652), .Y(n1859) );
  OAI21X1 U3558 ( .A(n6478), .B(n6649), .C(n1860), .Y(n4242) );
  NAND2X1 U3559 ( .A(\Mem[61][4] ), .B(n6653), .Y(n1860) );
  OAI21X1 U3560 ( .A(n6473), .B(n6649), .C(n1861), .Y(n4243) );
  NAND2X1 U3561 ( .A(\Mem[61][5] ), .B(n6652), .Y(n1861) );
  OAI21X1 U3562 ( .A(n6468), .B(n6649), .C(n1862), .Y(n4244) );
  NAND2X1 U3563 ( .A(\Mem[61][6] ), .B(n6652), .Y(n1862) );
  OAI21X1 U3564 ( .A(n6463), .B(n6649), .C(n1863), .Y(n4245) );
  NAND2X1 U3565 ( .A(\Mem[61][7] ), .B(n6652), .Y(n1863) );
  OAI21X1 U3566 ( .A(n6458), .B(n6649), .C(n1864), .Y(n4246) );
  NAND2X1 U3567 ( .A(\Mem[61][8] ), .B(n6652), .Y(n1864) );
  OAI21X1 U3568 ( .A(n6453), .B(n6649), .C(n1865), .Y(n4247) );
  NAND2X1 U3569 ( .A(\Mem[61][9] ), .B(n6652), .Y(n1865) );
  OAI21X1 U3570 ( .A(n6603), .B(n6649), .C(n1866), .Y(n4248) );
  NAND2X1 U3571 ( .A(\Mem[61][10] ), .B(n6652), .Y(n1866) );
  OAI21X1 U3572 ( .A(n6598), .B(n6649), .C(n1867), .Y(n4249) );
  NAND2X1 U3573 ( .A(\Mem[61][11] ), .B(n6652), .Y(n1867) );
  OAI21X1 U3574 ( .A(n6593), .B(n6649), .C(n1868), .Y(n4250) );
  NAND2X1 U3575 ( .A(\Mem[61][12] ), .B(n6652), .Y(n1868) );
  OAI21X1 U3576 ( .A(n6588), .B(n6650), .C(n1869), .Y(n4251) );
  NAND2X1 U3577 ( .A(\Mem[61][13] ), .B(n6652), .Y(n1869) );
  OAI21X1 U3578 ( .A(n6583), .B(n6650), .C(n1870), .Y(n4252) );
  NAND2X1 U3579 ( .A(\Mem[61][14] ), .B(n6652), .Y(n1870) );
  OAI21X1 U3580 ( .A(n6578), .B(n6650), .C(n1871), .Y(n4253) );
  NAND2X1 U3581 ( .A(\Mem[61][15] ), .B(n6651), .Y(n1871) );
  OAI21X1 U3582 ( .A(n6573), .B(n6650), .C(n1872), .Y(n4254) );
  NAND2X1 U3583 ( .A(\Mem[61][16] ), .B(n6652), .Y(n1872) );
  OAI21X1 U3584 ( .A(n6568), .B(n6650), .C(n1873), .Y(n4255) );
  NAND2X1 U3585 ( .A(\Mem[61][17] ), .B(n6651), .Y(n1873) );
  OAI21X1 U3586 ( .A(n6563), .B(n6650), .C(n1874), .Y(n4256) );
  NAND2X1 U3587 ( .A(\Mem[61][18] ), .B(n6651), .Y(n1874) );
  OAI21X1 U3588 ( .A(n6558), .B(n6650), .C(n1875), .Y(n4257) );
  NAND2X1 U3589 ( .A(\Mem[61][19] ), .B(n6651), .Y(n1875) );
  OAI21X1 U3590 ( .A(n6548), .B(n6650), .C(n1876), .Y(n4258) );
  NAND2X1 U3591 ( .A(\Mem[61][20] ), .B(n6651), .Y(n1876) );
  OAI21X1 U3592 ( .A(n6543), .B(n6650), .C(n1877), .Y(n4259) );
  NAND2X1 U3593 ( .A(\Mem[61][21] ), .B(n6651), .Y(n1877) );
  OAI21X1 U3594 ( .A(n6538), .B(n6650), .C(n1878), .Y(n4260) );
  NAND2X1 U3595 ( .A(\Mem[61][22] ), .B(n6652), .Y(n1878) );
  OAI21X1 U3596 ( .A(n6533), .B(n6651), .C(n1879), .Y(n4261) );
  NAND2X1 U3597 ( .A(\Mem[61][23] ), .B(n6651), .Y(n1879) );
  OAI21X1 U3598 ( .A(n6528), .B(n6650), .C(n1880), .Y(n4262) );
  NAND2X1 U3599 ( .A(\Mem[61][24] ), .B(n6652), .Y(n1880) );
  OAI21X1 U3600 ( .A(n6523), .B(n6651), .C(n1881), .Y(n4263) );
  NAND2X1 U3601 ( .A(\Mem[61][25] ), .B(n6652), .Y(n1881) );
  OAI21X1 U3602 ( .A(n6518), .B(n6651), .C(n1882), .Y(n4264) );
  NAND2X1 U3603 ( .A(\Mem[61][26] ), .B(n6652), .Y(n1882) );
  OAI21X1 U3604 ( .A(n6513), .B(n6651), .C(n1883), .Y(n4265) );
  NAND2X1 U3605 ( .A(\Mem[61][27] ), .B(n6652), .Y(n1883) );
  OAI21X1 U3606 ( .A(n6508), .B(n6651), .C(n1884), .Y(n4266) );
  NAND2X1 U3607 ( .A(\Mem[61][28] ), .B(n6652), .Y(n1884) );
  OAI21X1 U3608 ( .A(n6503), .B(n6651), .C(n1885), .Y(n4267) );
  NAND2X1 U3609 ( .A(\Mem[61][29] ), .B(n6652), .Y(n1885) );
  OAI21X1 U3610 ( .A(n6493), .B(n6651), .C(n1886), .Y(n4268) );
  NAND2X1 U3611 ( .A(\Mem[61][30] ), .B(n6653), .Y(n1886) );
  OAI21X1 U3612 ( .A(n6488), .B(n6651), .C(n1887), .Y(n4269) );
  NAND2X1 U3613 ( .A(\Mem[61][31] ), .B(n6653), .Y(n1887) );
  NAND2X1 U3614 ( .A(n7008), .B(n7023), .Y(n1855) );
  OAI21X1 U3615 ( .A(n6608), .B(n6645), .C(n1889), .Y(n4270) );
  NAND2X1 U3616 ( .A(\Mem[62][0] ), .B(n6648), .Y(n1889) );
  OAI21X1 U3617 ( .A(n6553), .B(n6644), .C(n1890), .Y(n4271) );
  NAND2X1 U3618 ( .A(\Mem[62][1] ), .B(n6648), .Y(n1890) );
  OAI21X1 U3619 ( .A(n6498), .B(n6644), .C(n1891), .Y(n4272) );
  NAND2X1 U3620 ( .A(\Mem[62][2] ), .B(n6648), .Y(n1891) );
  OAI21X1 U3621 ( .A(n6483), .B(n6644), .C(n1892), .Y(n4273) );
  NAND2X1 U3622 ( .A(\Mem[62][3] ), .B(n6647), .Y(n1892) );
  OAI21X1 U3623 ( .A(n6478), .B(n6644), .C(n1893), .Y(n4274) );
  NAND2X1 U3624 ( .A(\Mem[62][4] ), .B(n6648), .Y(n1893) );
  OAI21X1 U3625 ( .A(n6473), .B(n6644), .C(n1894), .Y(n4275) );
  NAND2X1 U3626 ( .A(\Mem[62][5] ), .B(n6647), .Y(n1894) );
  OAI21X1 U3627 ( .A(n6468), .B(n6644), .C(n1895), .Y(n4276) );
  NAND2X1 U3628 ( .A(\Mem[62][6] ), .B(n6647), .Y(n1895) );
  OAI21X1 U3629 ( .A(n6463), .B(n6644), .C(n1896), .Y(n4277) );
  NAND2X1 U3630 ( .A(\Mem[62][7] ), .B(n6647), .Y(n1896) );
  OAI21X1 U3631 ( .A(n6458), .B(n6644), .C(n1897), .Y(n4278) );
  NAND2X1 U3632 ( .A(\Mem[62][8] ), .B(n6647), .Y(n1897) );
  OAI21X1 U3633 ( .A(n6453), .B(n6644), .C(n1898), .Y(n4279) );
  NAND2X1 U3634 ( .A(\Mem[62][9] ), .B(n6647), .Y(n1898) );
  OAI21X1 U3635 ( .A(n6603), .B(n6644), .C(n1899), .Y(n4280) );
  NAND2X1 U3636 ( .A(\Mem[62][10] ), .B(n6647), .Y(n1899) );
  OAI21X1 U3637 ( .A(n6598), .B(n6644), .C(n1900), .Y(n4281) );
  NAND2X1 U3638 ( .A(\Mem[62][11] ), .B(n6647), .Y(n1900) );
  OAI21X1 U3639 ( .A(n6593), .B(n6644), .C(n1901), .Y(n4282) );
  NAND2X1 U3640 ( .A(\Mem[62][12] ), .B(n6647), .Y(n1901) );
  OAI21X1 U3641 ( .A(n6588), .B(n6645), .C(n1902), .Y(n4283) );
  NAND2X1 U3642 ( .A(\Mem[62][13] ), .B(n6647), .Y(n1902) );
  OAI21X1 U3643 ( .A(n6583), .B(n6645), .C(n1903), .Y(n4284) );
  NAND2X1 U3644 ( .A(\Mem[62][14] ), .B(n6647), .Y(n1903) );
  OAI21X1 U3645 ( .A(n6578), .B(n6645), .C(n1904), .Y(n4285) );
  NAND2X1 U3646 ( .A(\Mem[62][15] ), .B(n6646), .Y(n1904) );
  OAI21X1 U3647 ( .A(n6573), .B(n6645), .C(n1905), .Y(n4286) );
  NAND2X1 U3648 ( .A(\Mem[62][16] ), .B(n6647), .Y(n1905) );
  OAI21X1 U3649 ( .A(n6568), .B(n6645), .C(n1906), .Y(n4287) );
  NAND2X1 U3650 ( .A(\Mem[62][17] ), .B(n6646), .Y(n1906) );
  OAI21X1 U3651 ( .A(n6563), .B(n6645), .C(n1907), .Y(n4288) );
  NAND2X1 U3652 ( .A(\Mem[62][18] ), .B(n6646), .Y(n1907) );
  OAI21X1 U3653 ( .A(n6558), .B(n6645), .C(n1908), .Y(n4289) );
  NAND2X1 U3654 ( .A(\Mem[62][19] ), .B(n6646), .Y(n1908) );
  OAI21X1 U3655 ( .A(n6548), .B(n6645), .C(n1909), .Y(n4290) );
  NAND2X1 U3656 ( .A(\Mem[62][20] ), .B(n6646), .Y(n1909) );
  OAI21X1 U3657 ( .A(n6543), .B(n6645), .C(n1910), .Y(n4291) );
  NAND2X1 U3658 ( .A(\Mem[62][21] ), .B(n6646), .Y(n1910) );
  OAI21X1 U3659 ( .A(n6538), .B(n6645), .C(n1911), .Y(n4292) );
  NAND2X1 U3660 ( .A(\Mem[62][22] ), .B(n6647), .Y(n1911) );
  OAI21X1 U3661 ( .A(n6533), .B(n6646), .C(n1912), .Y(n4293) );
  NAND2X1 U3662 ( .A(\Mem[62][23] ), .B(n6646), .Y(n1912) );
  OAI21X1 U3663 ( .A(n6528), .B(n6645), .C(n1913), .Y(n4294) );
  NAND2X1 U3664 ( .A(\Mem[62][24] ), .B(n6647), .Y(n1913) );
  OAI21X1 U3665 ( .A(n6523), .B(n6646), .C(n1914), .Y(n4295) );
  NAND2X1 U3666 ( .A(\Mem[62][25] ), .B(n6647), .Y(n1914) );
  OAI21X1 U3667 ( .A(n6518), .B(n6646), .C(n1915), .Y(n4296) );
  NAND2X1 U3668 ( .A(\Mem[62][26] ), .B(n6647), .Y(n1915) );
  OAI21X1 U3669 ( .A(n6513), .B(n6646), .C(n1916), .Y(n4297) );
  NAND2X1 U3670 ( .A(\Mem[62][27] ), .B(n6647), .Y(n1916) );
  OAI21X1 U3671 ( .A(n6508), .B(n6646), .C(n1917), .Y(n4298) );
  NAND2X1 U3672 ( .A(\Mem[62][28] ), .B(n6647), .Y(n1917) );
  OAI21X1 U3673 ( .A(n6503), .B(n6646), .C(n1918), .Y(n4299) );
  NAND2X1 U3674 ( .A(\Mem[62][29] ), .B(n6647), .Y(n1918) );
  OAI21X1 U3675 ( .A(n6493), .B(n6646), .C(n1919), .Y(n4300) );
  NAND2X1 U3676 ( .A(\Mem[62][30] ), .B(n6648), .Y(n1919) );
  OAI21X1 U3677 ( .A(n6488), .B(n6646), .C(n1920), .Y(n4301) );
  NAND2X1 U3678 ( .A(\Mem[62][31] ), .B(n6648), .Y(n1920) );
  NAND2X1 U3679 ( .A(n7008), .B(n7024), .Y(n1888) );
  OAI21X1 U3680 ( .A(n6608), .B(n6640), .C(n1922), .Y(n4302) );
  NAND2X1 U3681 ( .A(\Mem[63][0] ), .B(n6643), .Y(n1922) );
  OAI21X1 U3682 ( .A(n6553), .B(n6639), .C(n1923), .Y(n4303) );
  NAND2X1 U3683 ( .A(\Mem[63][1] ), .B(n6643), .Y(n1923) );
  OAI21X1 U3684 ( .A(n6498), .B(n6639), .C(n1924), .Y(n4304) );
  NAND2X1 U3685 ( .A(\Mem[63][2] ), .B(n6643), .Y(n1924) );
  OAI21X1 U3686 ( .A(n6483), .B(n6639), .C(n1925), .Y(n4305) );
  NAND2X1 U3687 ( .A(\Mem[63][3] ), .B(n6642), .Y(n1925) );
  OAI21X1 U3688 ( .A(n6478), .B(n6639), .C(n1926), .Y(n4306) );
  NAND2X1 U3689 ( .A(\Mem[63][4] ), .B(n6643), .Y(n1926) );
  OAI21X1 U3690 ( .A(n6473), .B(n6639), .C(n1927), .Y(n4307) );
  NAND2X1 U3691 ( .A(\Mem[63][5] ), .B(n6642), .Y(n1927) );
  OAI21X1 U3692 ( .A(n6468), .B(n6639), .C(n1928), .Y(n4308) );
  NAND2X1 U3693 ( .A(\Mem[63][6] ), .B(n6642), .Y(n1928) );
  OAI21X1 U3694 ( .A(n6463), .B(n6639), .C(n1929), .Y(n4309) );
  NAND2X1 U3695 ( .A(\Mem[63][7] ), .B(n6642), .Y(n1929) );
  OAI21X1 U3696 ( .A(n6458), .B(n6639), .C(n1930), .Y(n4310) );
  NAND2X1 U3697 ( .A(\Mem[63][8] ), .B(n6642), .Y(n1930) );
  OAI21X1 U3698 ( .A(n6453), .B(n6639), .C(n1931), .Y(n4311) );
  NAND2X1 U3699 ( .A(\Mem[63][9] ), .B(n6642), .Y(n1931) );
  OAI21X1 U3700 ( .A(n6603), .B(n6639), .C(n1932), .Y(n4312) );
  NAND2X1 U3701 ( .A(\Mem[63][10] ), .B(n6642), .Y(n1932) );
  OAI21X1 U3702 ( .A(n6598), .B(n6639), .C(n1933), .Y(n4313) );
  NAND2X1 U3703 ( .A(\Mem[63][11] ), .B(n6642), .Y(n1933) );
  OAI21X1 U3704 ( .A(n6593), .B(n6639), .C(n1934), .Y(n4314) );
  NAND2X1 U3705 ( .A(\Mem[63][12] ), .B(n6642), .Y(n1934) );
  OAI21X1 U3706 ( .A(n6588), .B(n6640), .C(n1935), .Y(n4315) );
  NAND2X1 U3707 ( .A(\Mem[63][13] ), .B(n6642), .Y(n1935) );
  OAI21X1 U3708 ( .A(n6583), .B(n6640), .C(n1936), .Y(n4316) );
  NAND2X1 U3709 ( .A(\Mem[63][14] ), .B(n6642), .Y(n1936) );
  OAI21X1 U3710 ( .A(n6578), .B(n6640), .C(n1937), .Y(n4317) );
  NAND2X1 U3711 ( .A(\Mem[63][15] ), .B(n6641), .Y(n1937) );
  OAI21X1 U3712 ( .A(n6573), .B(n6640), .C(n1938), .Y(n4318) );
  NAND2X1 U3713 ( .A(\Mem[63][16] ), .B(n6642), .Y(n1938) );
  OAI21X1 U3714 ( .A(n6568), .B(n6640), .C(n1939), .Y(n4319) );
  NAND2X1 U3715 ( .A(\Mem[63][17] ), .B(n6641), .Y(n1939) );
  OAI21X1 U3716 ( .A(n6563), .B(n6640), .C(n1940), .Y(n4320) );
  NAND2X1 U3717 ( .A(\Mem[63][18] ), .B(n6641), .Y(n1940) );
  OAI21X1 U3718 ( .A(n6558), .B(n6640), .C(n1941), .Y(n4321) );
  NAND2X1 U3719 ( .A(\Mem[63][19] ), .B(n6641), .Y(n1941) );
  OAI21X1 U3720 ( .A(n6548), .B(n6640), .C(n1942), .Y(n4322) );
  NAND2X1 U3721 ( .A(\Mem[63][20] ), .B(n6641), .Y(n1942) );
  OAI21X1 U3722 ( .A(n6543), .B(n6640), .C(n1943), .Y(n4323) );
  NAND2X1 U3723 ( .A(\Mem[63][21] ), .B(n6641), .Y(n1943) );
  OAI21X1 U3724 ( .A(n6538), .B(n6640), .C(n1944), .Y(n4324) );
  NAND2X1 U3725 ( .A(\Mem[63][22] ), .B(n6642), .Y(n1944) );
  OAI21X1 U3726 ( .A(n6533), .B(n6641), .C(n1945), .Y(n4325) );
  NAND2X1 U3727 ( .A(\Mem[63][23] ), .B(n6641), .Y(n1945) );
  OAI21X1 U3728 ( .A(n6528), .B(n6640), .C(n1946), .Y(n4326) );
  NAND2X1 U3729 ( .A(\Mem[63][24] ), .B(n6642), .Y(n1946) );
  OAI21X1 U3730 ( .A(n6523), .B(n6641), .C(n1947), .Y(n4327) );
  NAND2X1 U3731 ( .A(\Mem[63][25] ), .B(n6642), .Y(n1947) );
  OAI21X1 U3732 ( .A(n6518), .B(n6641), .C(n1948), .Y(n4328) );
  NAND2X1 U3733 ( .A(\Mem[63][26] ), .B(n6642), .Y(n1948) );
  OAI21X1 U3734 ( .A(n6513), .B(n6641), .C(n1949), .Y(n4329) );
  NAND2X1 U3735 ( .A(\Mem[63][27] ), .B(n6642), .Y(n1949) );
  OAI21X1 U3736 ( .A(n6508), .B(n6641), .C(n1950), .Y(n4330) );
  NAND2X1 U3737 ( .A(\Mem[63][28] ), .B(n6642), .Y(n1950) );
  OAI21X1 U3738 ( .A(n6503), .B(n6641), .C(n1951), .Y(n4331) );
  NAND2X1 U3739 ( .A(\Mem[63][29] ), .B(n6642), .Y(n1951) );
  OAI21X1 U3740 ( .A(n6493), .B(n6641), .C(n1952), .Y(n4332) );
  NAND2X1 U3741 ( .A(\Mem[63][30] ), .B(n6643), .Y(n1952) );
  OAI21X1 U3742 ( .A(n6488), .B(n6641), .C(n1953), .Y(n4333) );
  NAND2X1 U3743 ( .A(\Mem[63][31] ), .B(n6643), .Y(n1953) );
  NAND2X1 U3744 ( .A(n7008), .B(n7021), .Y(n1921) );
  NAND3X1 U3746 ( .A(ADDR_WR[2]), .B(ADDR_WR[1]), .C(ADDR_WR[0]), .Y(n1954) );
  NAND3X1 U3748 ( .A(ADDR_WR[4]), .B(ADDR_WR[3]), .C(n80), .Y(n1955) );
  NOR2X1 U3749 ( .A(n7013), .B(n1957), .Y(n1156) );
  AOI22X1 U3752 ( .A(DOUT[0]), .B(n6938), .C(n6931), .D(N112), .Y(n1958) );
  AOI22X1 U3754 ( .A(DOUT[1]), .B(n6938), .C(N111), .D(n6931), .Y(n1960) );
  AOI22X1 U3756 ( .A(DOUT[2]), .B(n6937), .C(N110), .D(n6931), .Y(n1961) );
  AOI22X1 U3758 ( .A(DOUT[3]), .B(n6937), .C(N109), .D(n6931), .Y(n1962) );
  AOI22X1 U3760 ( .A(DOUT[4]), .B(n6937), .C(N108), .D(n6931), .Y(n1963) );
  AOI22X1 U3762 ( .A(DOUT[5]), .B(n6937), .C(N107), .D(n6931), .Y(n1964) );
  AOI22X1 U3764 ( .A(DOUT[6]), .B(n6937), .C(N106), .D(n6930), .Y(n1965) );
  AOI22X1 U3766 ( .A(DOUT[7]), .B(n6937), .C(N105), .D(n6930), .Y(n1966) );
  AOI22X1 U3768 ( .A(DOUT[8]), .B(n6937), .C(N104), .D(n6930), .Y(n1967) );
  AOI22X1 U3770 ( .A(DOUT[9]), .B(n6936), .C(N103), .D(n6930), .Y(n1968) );
  AOI22X1 U3772 ( .A(DOUT[10]), .B(n6936), .C(N102), .D(n6930), .Y(n1969) );
  AOI22X1 U3774 ( .A(DOUT[11]), .B(n6936), .C(N101), .D(n6930), .Y(n1970) );
  AOI22X1 U3776 ( .A(DOUT[12]), .B(n6936), .C(N100), .D(n6930), .Y(n1971) );
  AOI22X1 U3778 ( .A(DOUT[13]), .B(n6936), .C(N99), .D(n6930), .Y(n1972) );
  AOI22X1 U3780 ( .A(DOUT[14]), .B(n6936), .C(N98), .D(n6930), .Y(n1973) );
  AOI22X1 U3782 ( .A(DOUT[15]), .B(n6936), .C(N97), .D(n6930), .Y(n1974) );
  AOI22X1 U3784 ( .A(DOUT[16]), .B(n6935), .C(N96), .D(n6930), .Y(n1975) );
  AOI22X1 U3786 ( .A(DOUT[17]), .B(n6935), .C(N95), .D(n6930), .Y(n1976) );
  AOI22X1 U3788 ( .A(DOUT[18]), .B(n6935), .C(N94), .D(n6930), .Y(n1977) );
  AOI22X1 U3790 ( .A(DOUT[19]), .B(n6935), .C(N93), .D(n6929), .Y(n1978) );
  AOI22X1 U3792 ( .A(DOUT[20]), .B(n6935), .C(N92), .D(n6929), .Y(n1979) );
  AOI22X1 U3794 ( .A(DOUT[21]), .B(n6935), .C(N91), .D(n6929), .Y(n1980) );
  AOI22X1 U3796 ( .A(DOUT[22]), .B(n6935), .C(N90), .D(n6929), .Y(n1981) );
  AOI22X1 U3798 ( .A(DOUT[23]), .B(n6934), .C(N89), .D(n6929), .Y(n1982) );
  AOI22X1 U3800 ( .A(DOUT[24]), .B(n6934), .C(N88), .D(n6929), .Y(n1983) );
  AOI22X1 U3802 ( .A(DOUT[25]), .B(n6934), .C(N87), .D(n6929), .Y(n1984) );
  AOI22X1 U3804 ( .A(DOUT[26]), .B(n6933), .C(N86), .D(n6929), .Y(n1985) );
  AOI22X1 U3806 ( .A(DOUT[27]), .B(n6933), .C(N85), .D(n6929), .Y(n1986) );
  AOI22X1 U3808 ( .A(DOUT[28]), .B(n6933), .C(N84), .D(n6929), .Y(n1987) );
  AOI22X1 U3810 ( .A(DOUT[29]), .B(n6932), .C(N83), .D(n6929), .Y(n1988) );
  AOI22X1 U3812 ( .A(DOUT[30]), .B(n6932), .C(N82), .D(n6929), .Y(n1989) );
  AOI22X1 U3815 ( .A(DOUT[31]), .B(n6932), .C(N81), .D(n6929), .Y(n1990) );
  OAI21X1 U3817 ( .A(n6608), .B(n6635), .C(n1992), .Y(n2286) );
  NAND2X1 U3818 ( .A(\Mem[0][0] ), .B(n6638), .Y(n1992) );
  OAI21X1 U3819 ( .A(n6553), .B(n6634), .C(n1993), .Y(n2287) );
  NAND2X1 U3820 ( .A(\Mem[0][1] ), .B(n6638), .Y(n1993) );
  OAI21X1 U3821 ( .A(n6498), .B(n6634), .C(n1994), .Y(n2288) );
  NAND2X1 U3822 ( .A(\Mem[0][2] ), .B(n6638), .Y(n1994) );
  OAI21X1 U3823 ( .A(n6483), .B(n6634), .C(n1995), .Y(n2289) );
  NAND2X1 U3824 ( .A(\Mem[0][3] ), .B(n6637), .Y(n1995) );
  OAI21X1 U3825 ( .A(n6478), .B(n6634), .C(n1996), .Y(n2290) );
  NAND2X1 U3826 ( .A(\Mem[0][4] ), .B(n6638), .Y(n1996) );
  OAI21X1 U3827 ( .A(n6473), .B(n6634), .C(n1997), .Y(n2291) );
  NAND2X1 U3828 ( .A(\Mem[0][5] ), .B(n6637), .Y(n1997) );
  OAI21X1 U3829 ( .A(n6468), .B(n6634), .C(n1998), .Y(n2292) );
  NAND2X1 U3830 ( .A(\Mem[0][6] ), .B(n6637), .Y(n1998) );
  OAI21X1 U3831 ( .A(n6463), .B(n6634), .C(n1999), .Y(n2293) );
  NAND2X1 U3832 ( .A(\Mem[0][7] ), .B(n6637), .Y(n1999) );
  OAI21X1 U3833 ( .A(n6458), .B(n6634), .C(n2000), .Y(n2294) );
  NAND2X1 U3834 ( .A(\Mem[0][8] ), .B(n6637), .Y(n2000) );
  OAI21X1 U3835 ( .A(n6453), .B(n6634), .C(n2001), .Y(n2295) );
  NAND2X1 U3836 ( .A(\Mem[0][9] ), .B(n6637), .Y(n2001) );
  OAI21X1 U3837 ( .A(n6603), .B(n6634), .C(n2002), .Y(n2296) );
  NAND2X1 U3838 ( .A(\Mem[0][10] ), .B(n6637), .Y(n2002) );
  OAI21X1 U3839 ( .A(n6598), .B(n6634), .C(n2003), .Y(n2297) );
  NAND2X1 U3840 ( .A(\Mem[0][11] ), .B(n6637), .Y(n2003) );
  OAI21X1 U3841 ( .A(n6593), .B(n6634), .C(n2004), .Y(n2298) );
  NAND2X1 U3842 ( .A(\Mem[0][12] ), .B(n6637), .Y(n2004) );
  OAI21X1 U3843 ( .A(n6588), .B(n6635), .C(n2005), .Y(n2299) );
  NAND2X1 U3844 ( .A(\Mem[0][13] ), .B(n6637), .Y(n2005) );
  OAI21X1 U3845 ( .A(n6583), .B(n6635), .C(n2006), .Y(n2300) );
  NAND2X1 U3846 ( .A(\Mem[0][14] ), .B(n6637), .Y(n2006) );
  OAI21X1 U3847 ( .A(n6578), .B(n6635), .C(n2007), .Y(n2301) );
  NAND2X1 U3848 ( .A(\Mem[0][15] ), .B(n6636), .Y(n2007) );
  OAI21X1 U3849 ( .A(n6573), .B(n6635), .C(n2008), .Y(n2302) );
  NAND2X1 U3850 ( .A(\Mem[0][16] ), .B(n6637), .Y(n2008) );
  OAI21X1 U3851 ( .A(n6568), .B(n6635), .C(n2009), .Y(n2303) );
  NAND2X1 U3852 ( .A(\Mem[0][17] ), .B(n6636), .Y(n2009) );
  OAI21X1 U3853 ( .A(n6563), .B(n6635), .C(n2010), .Y(n2304) );
  NAND2X1 U3854 ( .A(\Mem[0][18] ), .B(n6636), .Y(n2010) );
  OAI21X1 U3855 ( .A(n6558), .B(n6635), .C(n2011), .Y(n2305) );
  NAND2X1 U3856 ( .A(\Mem[0][19] ), .B(n6636), .Y(n2011) );
  OAI21X1 U3857 ( .A(n6548), .B(n6635), .C(n2012), .Y(n2306) );
  NAND2X1 U3858 ( .A(\Mem[0][20] ), .B(n6636), .Y(n2012) );
  OAI21X1 U3859 ( .A(n6543), .B(n6635), .C(n2013), .Y(n2307) );
  NAND2X1 U3860 ( .A(\Mem[0][21] ), .B(n6636), .Y(n2013) );
  OAI21X1 U3861 ( .A(n6538), .B(n6635), .C(n2014), .Y(n2308) );
  NAND2X1 U3862 ( .A(\Mem[0][22] ), .B(n6637), .Y(n2014) );
  OAI21X1 U3863 ( .A(n6533), .B(n6636), .C(n2015), .Y(n2309) );
  NAND2X1 U3864 ( .A(\Mem[0][23] ), .B(n6636), .Y(n2015) );
  OAI21X1 U3865 ( .A(n6528), .B(n6635), .C(n2016), .Y(n2310) );
  NAND2X1 U3866 ( .A(\Mem[0][24] ), .B(n6637), .Y(n2016) );
  OAI21X1 U3867 ( .A(n6523), .B(n6636), .C(n2017), .Y(n2311) );
  NAND2X1 U3868 ( .A(\Mem[0][25] ), .B(n6637), .Y(n2017) );
  OAI21X1 U3869 ( .A(n6518), .B(n6636), .C(n2018), .Y(n2312) );
  NAND2X1 U3870 ( .A(\Mem[0][26] ), .B(n6637), .Y(n2018) );
  OAI21X1 U3871 ( .A(n6513), .B(n6636), .C(n2019), .Y(n2313) );
  NAND2X1 U3872 ( .A(\Mem[0][27] ), .B(n6637), .Y(n2019) );
  OAI21X1 U3873 ( .A(n6508), .B(n6636), .C(n2020), .Y(n2314) );
  NAND2X1 U3874 ( .A(\Mem[0][28] ), .B(n6637), .Y(n2020) );
  OAI21X1 U3875 ( .A(n6503), .B(n6636), .C(n2021), .Y(n2315) );
  NAND2X1 U3876 ( .A(\Mem[0][29] ), .B(n6637), .Y(n2021) );
  OAI21X1 U3877 ( .A(n6493), .B(n6636), .C(n2022), .Y(n2316) );
  NAND2X1 U3878 ( .A(\Mem[0][30] ), .B(n6638), .Y(n2022) );
  OAI21X1 U3879 ( .A(n6488), .B(n6636), .C(n2023), .Y(n2317) );
  NAND2X1 U3880 ( .A(\Mem[0][31] ), .B(n6638), .Y(n2023) );
  NAND2X1 U3881 ( .A(n7016), .B(n7004), .Y(n1991) );
  NAND3X1 U3883 ( .A(n7025), .B(n7020), .C(n7026), .Y(n2024) );
  OAI21X1 U3884 ( .A(n6608), .B(n6630), .C(n2029), .Y(n2318) );
  NAND2X1 U3885 ( .A(\Mem[1][0] ), .B(n6633), .Y(n2029) );
  OAI21X1 U3886 ( .A(n6553), .B(n6629), .C(n2030), .Y(n2319) );
  NAND2X1 U3887 ( .A(\Mem[1][1] ), .B(n6633), .Y(n2030) );
  OAI21X1 U3888 ( .A(n6498), .B(n6629), .C(n2031), .Y(n2320) );
  NAND2X1 U3889 ( .A(\Mem[1][2] ), .B(n6633), .Y(n2031) );
  OAI21X1 U3890 ( .A(n6483), .B(n6629), .C(n2032), .Y(n2321) );
  NAND2X1 U3891 ( .A(\Mem[1][3] ), .B(n6632), .Y(n2032) );
  OAI21X1 U3892 ( .A(n6478), .B(n6629), .C(n2033), .Y(n2322) );
  NAND2X1 U3893 ( .A(\Mem[1][4] ), .B(n6633), .Y(n2033) );
  OAI21X1 U3894 ( .A(n6473), .B(n6629), .C(n2034), .Y(n2323) );
  NAND2X1 U3895 ( .A(\Mem[1][5] ), .B(n6632), .Y(n2034) );
  OAI21X1 U3896 ( .A(n6468), .B(n6629), .C(n2035), .Y(n2324) );
  NAND2X1 U3897 ( .A(\Mem[1][6] ), .B(n6632), .Y(n2035) );
  OAI21X1 U3898 ( .A(n6463), .B(n6629), .C(n2036), .Y(n2325) );
  NAND2X1 U3899 ( .A(\Mem[1][7] ), .B(n6632), .Y(n2036) );
  OAI21X1 U3900 ( .A(n6458), .B(n6629), .C(n2037), .Y(n2326) );
  NAND2X1 U3901 ( .A(\Mem[1][8] ), .B(n6632), .Y(n2037) );
  OAI21X1 U3902 ( .A(n6453), .B(n6629), .C(n2038), .Y(n2327) );
  NAND2X1 U3903 ( .A(\Mem[1][9] ), .B(n6632), .Y(n2038) );
  OAI21X1 U3904 ( .A(n6603), .B(n6629), .C(n2039), .Y(n2328) );
  NAND2X1 U3905 ( .A(\Mem[1][10] ), .B(n6632), .Y(n2039) );
  OAI21X1 U3906 ( .A(n6598), .B(n6629), .C(n2040), .Y(n2329) );
  NAND2X1 U3907 ( .A(\Mem[1][11] ), .B(n6632), .Y(n2040) );
  OAI21X1 U3908 ( .A(n6593), .B(n6629), .C(n2041), .Y(n2330) );
  NAND2X1 U3909 ( .A(\Mem[1][12] ), .B(n6632), .Y(n2041) );
  OAI21X1 U3910 ( .A(n6588), .B(n6630), .C(n2042), .Y(n2331) );
  NAND2X1 U3911 ( .A(\Mem[1][13] ), .B(n6632), .Y(n2042) );
  OAI21X1 U3912 ( .A(n6583), .B(n6630), .C(n2043), .Y(n2332) );
  NAND2X1 U3913 ( .A(\Mem[1][14] ), .B(n6632), .Y(n2043) );
  OAI21X1 U3914 ( .A(n6578), .B(n6630), .C(n2044), .Y(n2333) );
  NAND2X1 U3915 ( .A(\Mem[1][15] ), .B(n6631), .Y(n2044) );
  OAI21X1 U3916 ( .A(n6573), .B(n6630), .C(n2045), .Y(n2334) );
  NAND2X1 U3917 ( .A(\Mem[1][16] ), .B(n6632), .Y(n2045) );
  OAI21X1 U3918 ( .A(n6568), .B(n6630), .C(n2046), .Y(n2335) );
  NAND2X1 U3919 ( .A(\Mem[1][17] ), .B(n6631), .Y(n2046) );
  OAI21X1 U3920 ( .A(n6563), .B(n6630), .C(n2047), .Y(n2336) );
  NAND2X1 U3921 ( .A(\Mem[1][18] ), .B(n6631), .Y(n2047) );
  OAI21X1 U3922 ( .A(n6558), .B(n6630), .C(n2048), .Y(n2337) );
  NAND2X1 U3923 ( .A(\Mem[1][19] ), .B(n6631), .Y(n2048) );
  OAI21X1 U3924 ( .A(n6548), .B(n6630), .C(n2049), .Y(n2338) );
  NAND2X1 U3925 ( .A(\Mem[1][20] ), .B(n6631), .Y(n2049) );
  OAI21X1 U3926 ( .A(n6543), .B(n6630), .C(n2050), .Y(n2339) );
  NAND2X1 U3927 ( .A(\Mem[1][21] ), .B(n6631), .Y(n2050) );
  OAI21X1 U3928 ( .A(n6538), .B(n6630), .C(n2051), .Y(n2340) );
  NAND2X1 U3929 ( .A(\Mem[1][22] ), .B(n6632), .Y(n2051) );
  OAI21X1 U3930 ( .A(n6533), .B(n6631), .C(n2052), .Y(n2341) );
  NAND2X1 U3931 ( .A(\Mem[1][23] ), .B(n6631), .Y(n2052) );
  OAI21X1 U3932 ( .A(n6528), .B(n6630), .C(n2053), .Y(n2342) );
  NAND2X1 U3933 ( .A(\Mem[1][24] ), .B(n6632), .Y(n2053) );
  OAI21X1 U3934 ( .A(n6523), .B(n6631), .C(n2054), .Y(n2343) );
  NAND2X1 U3935 ( .A(\Mem[1][25] ), .B(n6632), .Y(n2054) );
  OAI21X1 U3936 ( .A(n6518), .B(n6631), .C(n2055), .Y(n2344) );
  NAND2X1 U3937 ( .A(\Mem[1][26] ), .B(n6632), .Y(n2055) );
  OAI21X1 U3938 ( .A(n6513), .B(n6631), .C(n2056), .Y(n2345) );
  NAND2X1 U3939 ( .A(\Mem[1][27] ), .B(n6632), .Y(n2056) );
  OAI21X1 U3940 ( .A(n6508), .B(n6631), .C(n2057), .Y(n2346) );
  NAND2X1 U3941 ( .A(\Mem[1][28] ), .B(n6632), .Y(n2057) );
  OAI21X1 U3942 ( .A(n6503), .B(n6631), .C(n2058), .Y(n2347) );
  NAND2X1 U3943 ( .A(\Mem[1][29] ), .B(n6632), .Y(n2058) );
  OAI21X1 U3944 ( .A(n6493), .B(n6631), .C(n2059), .Y(n2348) );
  NAND2X1 U3945 ( .A(\Mem[1][30] ), .B(n6633), .Y(n2059) );
  OAI21X1 U3946 ( .A(n6488), .B(n6631), .C(n2060), .Y(n2349) );
  NAND2X1 U3947 ( .A(\Mem[1][31] ), .B(n6633), .Y(n2060) );
  NAND2X1 U3948 ( .A(n7017), .B(n7004), .Y(n2028) );
  NAND3X1 U3950 ( .A(n7025), .B(n7020), .C(ADDR_WR[0]), .Y(n2061) );
  OAI21X1 U3951 ( .A(n6608), .B(n6625), .C(n2063), .Y(n2350) );
  NAND2X1 U3952 ( .A(\Mem[2][0] ), .B(n6628), .Y(n2063) );
  OAI21X1 U3953 ( .A(n6553), .B(n6624), .C(n2064), .Y(n2351) );
  NAND2X1 U3954 ( .A(\Mem[2][1] ), .B(n6628), .Y(n2064) );
  OAI21X1 U3955 ( .A(n6498), .B(n6624), .C(n2065), .Y(n2352) );
  NAND2X1 U3956 ( .A(\Mem[2][2] ), .B(n6628), .Y(n2065) );
  OAI21X1 U3957 ( .A(n6483), .B(n6624), .C(n2066), .Y(n2353) );
  NAND2X1 U3958 ( .A(\Mem[2][3] ), .B(n6627), .Y(n2066) );
  OAI21X1 U3959 ( .A(n6478), .B(n6624), .C(n2067), .Y(n2354) );
  NAND2X1 U3960 ( .A(\Mem[2][4] ), .B(n6628), .Y(n2067) );
  OAI21X1 U3961 ( .A(n6473), .B(n6624), .C(n2068), .Y(n2355) );
  NAND2X1 U3962 ( .A(\Mem[2][5] ), .B(n6627), .Y(n2068) );
  OAI21X1 U3963 ( .A(n6468), .B(n6624), .C(n2069), .Y(n2356) );
  NAND2X1 U3964 ( .A(\Mem[2][6] ), .B(n6627), .Y(n2069) );
  OAI21X1 U3965 ( .A(n6463), .B(n6624), .C(n2070), .Y(n2357) );
  NAND2X1 U3966 ( .A(\Mem[2][7] ), .B(n6627), .Y(n2070) );
  OAI21X1 U3967 ( .A(n6458), .B(n6624), .C(n2071), .Y(n2358) );
  NAND2X1 U3968 ( .A(\Mem[2][8] ), .B(n6627), .Y(n2071) );
  OAI21X1 U3969 ( .A(n6453), .B(n6624), .C(n2072), .Y(n2359) );
  NAND2X1 U3970 ( .A(\Mem[2][9] ), .B(n6627), .Y(n2072) );
  OAI21X1 U3971 ( .A(n6603), .B(n6624), .C(n2073), .Y(n2360) );
  NAND2X1 U3972 ( .A(\Mem[2][10] ), .B(n6627), .Y(n2073) );
  OAI21X1 U3973 ( .A(n6598), .B(n6624), .C(n2074), .Y(n2361) );
  NAND2X1 U3974 ( .A(\Mem[2][11] ), .B(n6627), .Y(n2074) );
  OAI21X1 U3975 ( .A(n6593), .B(n6624), .C(n2075), .Y(n2362) );
  NAND2X1 U3976 ( .A(\Mem[2][12] ), .B(n6627), .Y(n2075) );
  OAI21X1 U3977 ( .A(n6588), .B(n6625), .C(n2076), .Y(n2363) );
  NAND2X1 U3978 ( .A(\Mem[2][13] ), .B(n6627), .Y(n2076) );
  OAI21X1 U3979 ( .A(n6583), .B(n6625), .C(n2077), .Y(n2364) );
  NAND2X1 U3980 ( .A(\Mem[2][14] ), .B(n6627), .Y(n2077) );
  OAI21X1 U3981 ( .A(n6578), .B(n6625), .C(n2078), .Y(n2365) );
  NAND2X1 U3982 ( .A(\Mem[2][15] ), .B(n6626), .Y(n2078) );
  OAI21X1 U3983 ( .A(n6573), .B(n6625), .C(n2079), .Y(n2366) );
  NAND2X1 U3984 ( .A(\Mem[2][16] ), .B(n6627), .Y(n2079) );
  OAI21X1 U3985 ( .A(n6568), .B(n6625), .C(n2080), .Y(n2367) );
  NAND2X1 U3986 ( .A(\Mem[2][17] ), .B(n6626), .Y(n2080) );
  OAI21X1 U3987 ( .A(n6563), .B(n6625), .C(n2081), .Y(n2368) );
  NAND2X1 U3988 ( .A(\Mem[2][18] ), .B(n6626), .Y(n2081) );
  OAI21X1 U3989 ( .A(n6558), .B(n6625), .C(n2082), .Y(n2369) );
  NAND2X1 U3990 ( .A(\Mem[2][19] ), .B(n6626), .Y(n2082) );
  OAI21X1 U3991 ( .A(n6548), .B(n6625), .C(n2083), .Y(n2370) );
  NAND2X1 U3992 ( .A(\Mem[2][20] ), .B(n6626), .Y(n2083) );
  OAI21X1 U3993 ( .A(n6543), .B(n6625), .C(n2084), .Y(n2371) );
  NAND2X1 U3994 ( .A(\Mem[2][21] ), .B(n6626), .Y(n2084) );
  OAI21X1 U3995 ( .A(n6538), .B(n6625), .C(n2085), .Y(n2372) );
  NAND2X1 U3996 ( .A(\Mem[2][22] ), .B(n6627), .Y(n2085) );
  OAI21X1 U3997 ( .A(n6533), .B(n6626), .C(n2086), .Y(n2373) );
  NAND2X1 U3998 ( .A(\Mem[2][23] ), .B(n6626), .Y(n2086) );
  OAI21X1 U3999 ( .A(n6528), .B(n6625), .C(n2087), .Y(n2374) );
  NAND2X1 U4000 ( .A(\Mem[2][24] ), .B(n6627), .Y(n2087) );
  OAI21X1 U4001 ( .A(n6523), .B(n6626), .C(n2088), .Y(n2375) );
  NAND2X1 U4002 ( .A(\Mem[2][25] ), .B(n6627), .Y(n2088) );
  OAI21X1 U4003 ( .A(n6518), .B(n6626), .C(n2089), .Y(n2376) );
  NAND2X1 U4004 ( .A(\Mem[2][26] ), .B(n6627), .Y(n2089) );
  OAI21X1 U4005 ( .A(n6513), .B(n6626), .C(n2090), .Y(n2377) );
  NAND2X1 U4006 ( .A(\Mem[2][27] ), .B(n6627), .Y(n2090) );
  OAI21X1 U4007 ( .A(n6508), .B(n6626), .C(n2091), .Y(n2378) );
  NAND2X1 U4008 ( .A(\Mem[2][28] ), .B(n6627), .Y(n2091) );
  OAI21X1 U4009 ( .A(n6503), .B(n6626), .C(n2092), .Y(n2379) );
  NAND2X1 U4010 ( .A(\Mem[2][29] ), .B(n6627), .Y(n2092) );
  OAI21X1 U4011 ( .A(n6493), .B(n6626), .C(n2093), .Y(n2380) );
  NAND2X1 U4012 ( .A(\Mem[2][30] ), .B(n6628), .Y(n2093) );
  OAI21X1 U4013 ( .A(n6488), .B(n6626), .C(n2094), .Y(n2381) );
  NAND2X1 U4014 ( .A(\Mem[2][31] ), .B(n6628), .Y(n2094) );
  NAND2X1 U4015 ( .A(n7018), .B(n7004), .Y(n2062) );
  NAND3X1 U4017 ( .A(n7026), .B(n7020), .C(ADDR_WR[1]), .Y(n2095) );
  OAI21X1 U4018 ( .A(n6608), .B(n6620), .C(n2097), .Y(n2382) );
  NAND2X1 U4019 ( .A(\Mem[3][0] ), .B(n6623), .Y(n2097) );
  OAI21X1 U4020 ( .A(n6553), .B(n6619), .C(n2098), .Y(n2383) );
  NAND2X1 U4021 ( .A(\Mem[3][1] ), .B(n6623), .Y(n2098) );
  OAI21X1 U4022 ( .A(n6498), .B(n6619), .C(n2099), .Y(n2384) );
  NAND2X1 U4023 ( .A(\Mem[3][2] ), .B(n6623), .Y(n2099) );
  OAI21X1 U4024 ( .A(n6483), .B(n6619), .C(n2100), .Y(n2385) );
  NAND2X1 U4025 ( .A(\Mem[3][3] ), .B(n6622), .Y(n2100) );
  OAI21X1 U4026 ( .A(n6478), .B(n6619), .C(n2101), .Y(n2386) );
  NAND2X1 U4027 ( .A(\Mem[3][4] ), .B(n6623), .Y(n2101) );
  OAI21X1 U4028 ( .A(n6473), .B(n6619), .C(n2102), .Y(n2387) );
  NAND2X1 U4029 ( .A(\Mem[3][5] ), .B(n6622), .Y(n2102) );
  OAI21X1 U4030 ( .A(n6468), .B(n6619), .C(n2103), .Y(n2388) );
  NAND2X1 U4031 ( .A(\Mem[3][6] ), .B(n6622), .Y(n2103) );
  OAI21X1 U4032 ( .A(n6463), .B(n6619), .C(n2104), .Y(n2389) );
  NAND2X1 U4033 ( .A(\Mem[3][7] ), .B(n6622), .Y(n2104) );
  OAI21X1 U4034 ( .A(n6458), .B(n6619), .C(n2105), .Y(n2390) );
  NAND2X1 U4035 ( .A(\Mem[3][8] ), .B(n6622), .Y(n2105) );
  OAI21X1 U4036 ( .A(n6453), .B(n6619), .C(n2106), .Y(n2391) );
  NAND2X1 U4037 ( .A(\Mem[3][9] ), .B(n6622), .Y(n2106) );
  OAI21X1 U4038 ( .A(n6603), .B(n6619), .C(n2107), .Y(n2392) );
  NAND2X1 U4039 ( .A(\Mem[3][10] ), .B(n6622), .Y(n2107) );
  OAI21X1 U4040 ( .A(n6598), .B(n6619), .C(n2108), .Y(n2393) );
  NAND2X1 U4041 ( .A(\Mem[3][11] ), .B(n6622), .Y(n2108) );
  OAI21X1 U4042 ( .A(n6593), .B(n6619), .C(n2109), .Y(n2394) );
  NAND2X1 U4043 ( .A(\Mem[3][12] ), .B(n6622), .Y(n2109) );
  OAI21X1 U4044 ( .A(n6588), .B(n6620), .C(n2110), .Y(n2395) );
  NAND2X1 U4045 ( .A(\Mem[3][13] ), .B(n6622), .Y(n2110) );
  OAI21X1 U4046 ( .A(n6583), .B(n6620), .C(n2111), .Y(n2396) );
  NAND2X1 U4047 ( .A(\Mem[3][14] ), .B(n6622), .Y(n2111) );
  OAI21X1 U4048 ( .A(n6578), .B(n6620), .C(n2112), .Y(n2397) );
  NAND2X1 U4049 ( .A(\Mem[3][15] ), .B(n6621), .Y(n2112) );
  OAI21X1 U4050 ( .A(n6573), .B(n6620), .C(n2113), .Y(n2398) );
  NAND2X1 U4051 ( .A(\Mem[3][16] ), .B(n6622), .Y(n2113) );
  OAI21X1 U4052 ( .A(n6568), .B(n6620), .C(n2114), .Y(n2399) );
  NAND2X1 U4053 ( .A(\Mem[3][17] ), .B(n6621), .Y(n2114) );
  OAI21X1 U4054 ( .A(n6563), .B(n6620), .C(n2115), .Y(n2400) );
  NAND2X1 U4055 ( .A(\Mem[3][18] ), .B(n6621), .Y(n2115) );
  OAI21X1 U4056 ( .A(n6558), .B(n6620), .C(n2116), .Y(n2401) );
  NAND2X1 U4057 ( .A(\Mem[3][19] ), .B(n6621), .Y(n2116) );
  OAI21X1 U4058 ( .A(n6548), .B(n6620), .C(n2117), .Y(n2402) );
  NAND2X1 U4059 ( .A(\Mem[3][20] ), .B(n6621), .Y(n2117) );
  OAI21X1 U4060 ( .A(n6543), .B(n6620), .C(n2118), .Y(n2403) );
  NAND2X1 U4061 ( .A(\Mem[3][21] ), .B(n6621), .Y(n2118) );
  OAI21X1 U4062 ( .A(n6538), .B(n6620), .C(n2119), .Y(n2404) );
  NAND2X1 U4063 ( .A(\Mem[3][22] ), .B(n6622), .Y(n2119) );
  OAI21X1 U4064 ( .A(n6533), .B(n6621), .C(n2120), .Y(n2405) );
  NAND2X1 U4065 ( .A(\Mem[3][23] ), .B(n6621), .Y(n2120) );
  OAI21X1 U4066 ( .A(n6528), .B(n6620), .C(n2121), .Y(n2406) );
  NAND2X1 U4067 ( .A(\Mem[3][24] ), .B(n6622), .Y(n2121) );
  OAI21X1 U4068 ( .A(n6523), .B(n6621), .C(n2122), .Y(n2407) );
  NAND2X1 U4069 ( .A(\Mem[3][25] ), .B(n6622), .Y(n2122) );
  OAI21X1 U4070 ( .A(n6518), .B(n6621), .C(n2123), .Y(n2408) );
  NAND2X1 U4071 ( .A(\Mem[3][26] ), .B(n6622), .Y(n2123) );
  OAI21X1 U4072 ( .A(n6513), .B(n6621), .C(n2124), .Y(n2409) );
  NAND2X1 U4073 ( .A(\Mem[3][27] ), .B(n6622), .Y(n2124) );
  OAI21X1 U4074 ( .A(n6508), .B(n6621), .C(n2125), .Y(n2410) );
  NAND2X1 U4075 ( .A(\Mem[3][28] ), .B(n6622), .Y(n2125) );
  OAI21X1 U4076 ( .A(n6503), .B(n6621), .C(n2126), .Y(n2411) );
  NAND2X1 U4077 ( .A(\Mem[3][29] ), .B(n6622), .Y(n2126) );
  OAI21X1 U4078 ( .A(n6493), .B(n6621), .C(n2127), .Y(n2412) );
  NAND2X1 U4079 ( .A(\Mem[3][30] ), .B(n6623), .Y(n2127) );
  OAI21X1 U4080 ( .A(n6488), .B(n6621), .C(n2128), .Y(n2413) );
  NAND2X1 U4081 ( .A(\Mem[3][31] ), .B(n6623), .Y(n2128) );
  NAND2X1 U4082 ( .A(n7019), .B(n7004), .Y(n2096) );
  NAND3X1 U4084 ( .A(ADDR_WR[1]), .B(n7020), .C(ADDR_WR[0]), .Y(n2129) );
  OAI21X1 U4086 ( .A(n6608), .B(n6615), .C(n2131), .Y(n2414) );
  NAND2X1 U4087 ( .A(\Mem[4][0] ), .B(n6618), .Y(n2131) );
  OAI21X1 U4088 ( .A(n6553), .B(n6614), .C(n2132), .Y(n2415) );
  NAND2X1 U4089 ( .A(\Mem[4][1] ), .B(n6618), .Y(n2132) );
  OAI21X1 U4090 ( .A(n6498), .B(n6614), .C(n2133), .Y(n2416) );
  NAND2X1 U4091 ( .A(\Mem[4][2] ), .B(n6618), .Y(n2133) );
  OAI21X1 U4092 ( .A(n6483), .B(n6614), .C(n2134), .Y(n2417) );
  NAND2X1 U4093 ( .A(\Mem[4][3] ), .B(n6617), .Y(n2134) );
  OAI21X1 U4094 ( .A(n6478), .B(n6614), .C(n2135), .Y(n2418) );
  NAND2X1 U4095 ( .A(\Mem[4][4] ), .B(n6618), .Y(n2135) );
  OAI21X1 U4096 ( .A(n6473), .B(n6614), .C(n2136), .Y(n2419) );
  NAND2X1 U4097 ( .A(\Mem[4][5] ), .B(n6617), .Y(n2136) );
  OAI21X1 U4098 ( .A(n6468), .B(n6614), .C(n2137), .Y(n2420) );
  NAND2X1 U4099 ( .A(\Mem[4][6] ), .B(n6617), .Y(n2137) );
  OAI21X1 U4100 ( .A(n6463), .B(n6614), .C(n2138), .Y(n2421) );
  NAND2X1 U4101 ( .A(\Mem[4][7] ), .B(n6617), .Y(n2138) );
  OAI21X1 U4102 ( .A(n6458), .B(n6614), .C(n2139), .Y(n2422) );
  NAND2X1 U4103 ( .A(\Mem[4][8] ), .B(n6617), .Y(n2139) );
  OAI21X1 U4104 ( .A(n6453), .B(n6614), .C(n2140), .Y(n2423) );
  NAND2X1 U4105 ( .A(\Mem[4][9] ), .B(n6617), .Y(n2140) );
  OAI21X1 U4106 ( .A(n6603), .B(n6614), .C(n2141), .Y(n2424) );
  NAND2X1 U4107 ( .A(\Mem[4][10] ), .B(n6617), .Y(n2141) );
  OAI21X1 U4108 ( .A(n6598), .B(n6614), .C(n2142), .Y(n2425) );
  NAND2X1 U4109 ( .A(\Mem[4][11] ), .B(n6617), .Y(n2142) );
  OAI21X1 U4110 ( .A(n6593), .B(n6614), .C(n2143), .Y(n2426) );
  NAND2X1 U4111 ( .A(\Mem[4][12] ), .B(n6617), .Y(n2143) );
  OAI21X1 U4112 ( .A(n6588), .B(n6615), .C(n2144), .Y(n2427) );
  NAND2X1 U4113 ( .A(\Mem[4][13] ), .B(n6617), .Y(n2144) );
  OAI21X1 U4114 ( .A(n6583), .B(n6615), .C(n2145), .Y(n2428) );
  NAND2X1 U4115 ( .A(\Mem[4][14] ), .B(n6617), .Y(n2145) );
  OAI21X1 U4116 ( .A(n6578), .B(n6615), .C(n2146), .Y(n2429) );
  NAND2X1 U4117 ( .A(\Mem[4][15] ), .B(n6616), .Y(n2146) );
  OAI21X1 U4118 ( .A(n6573), .B(n6615), .C(n2147), .Y(n2430) );
  NAND2X1 U4119 ( .A(\Mem[4][16] ), .B(n6617), .Y(n2147) );
  OAI21X1 U4120 ( .A(n6568), .B(n6615), .C(n2148), .Y(n2431) );
  NAND2X1 U4121 ( .A(\Mem[4][17] ), .B(n6616), .Y(n2148) );
  OAI21X1 U4122 ( .A(n6563), .B(n6615), .C(n2149), .Y(n2432) );
  NAND2X1 U4123 ( .A(\Mem[4][18] ), .B(n6616), .Y(n2149) );
  OAI21X1 U4124 ( .A(n6558), .B(n6615), .C(n2150), .Y(n2433) );
  NAND2X1 U4125 ( .A(\Mem[4][19] ), .B(n6616), .Y(n2150) );
  OAI21X1 U4126 ( .A(n6548), .B(n6615), .C(n2151), .Y(n2434) );
  NAND2X1 U4127 ( .A(\Mem[4][20] ), .B(n6616), .Y(n2151) );
  OAI21X1 U4128 ( .A(n6543), .B(n6615), .C(n2152), .Y(n2435) );
  NAND2X1 U4129 ( .A(\Mem[4][21] ), .B(n6616), .Y(n2152) );
  OAI21X1 U4130 ( .A(n6538), .B(n6615), .C(n2153), .Y(n2436) );
  NAND2X1 U4131 ( .A(\Mem[4][22] ), .B(n6617), .Y(n2153) );
  OAI21X1 U4132 ( .A(n6533), .B(n6616), .C(n2154), .Y(n2437) );
  NAND2X1 U4133 ( .A(\Mem[4][23] ), .B(n6616), .Y(n2154) );
  OAI21X1 U4134 ( .A(n6528), .B(n6615), .C(n2155), .Y(n2438) );
  NAND2X1 U4135 ( .A(\Mem[4][24] ), .B(n6617), .Y(n2155) );
  OAI21X1 U4136 ( .A(n6523), .B(n6616), .C(n2156), .Y(n2439) );
  NAND2X1 U4137 ( .A(\Mem[4][25] ), .B(n6617), .Y(n2156) );
  OAI21X1 U4138 ( .A(n6518), .B(n6616), .C(n2157), .Y(n2440) );
  NAND2X1 U4139 ( .A(\Mem[4][26] ), .B(n6617), .Y(n2157) );
  OAI21X1 U4140 ( .A(n6513), .B(n6616), .C(n2158), .Y(n2441) );
  NAND2X1 U4141 ( .A(\Mem[4][27] ), .B(n6617), .Y(n2158) );
  OAI21X1 U4142 ( .A(n6508), .B(n6616), .C(n2159), .Y(n2442) );
  NAND2X1 U4143 ( .A(\Mem[4][28] ), .B(n6617), .Y(n2159) );
  OAI21X1 U4144 ( .A(n6503), .B(n6616), .C(n2160), .Y(n2443) );
  NAND2X1 U4145 ( .A(\Mem[4][29] ), .B(n6617), .Y(n2160) );
  OAI21X1 U4146 ( .A(n6493), .B(n6616), .C(n2161), .Y(n2444) );
  NAND2X1 U4147 ( .A(\Mem[4][30] ), .B(n6618), .Y(n2161) );
  OAI21X1 U4148 ( .A(n6488), .B(n6616), .C(n2162), .Y(n2445) );
  NAND2X1 U4149 ( .A(\Mem[4][31] ), .B(n6618), .Y(n2162) );
  NAND2X1 U4150 ( .A(n7022), .B(n7004), .Y(n2130) );
  NAND3X1 U4152 ( .A(n7026), .B(n7025), .C(ADDR_WR[2]), .Y(n2163) );
  OAI21X1 U4153 ( .A(n6604), .B(n6610), .C(n2165), .Y(n2446) );
  NAND2X1 U4154 ( .A(\Mem[5][0] ), .B(n6613), .Y(n2165) );
  OAI21X1 U4155 ( .A(n6549), .B(n6609), .C(n2166), .Y(n2447) );
  NAND2X1 U4156 ( .A(\Mem[5][1] ), .B(n6613), .Y(n2166) );
  OAI21X1 U4157 ( .A(n6494), .B(n6609), .C(n2167), .Y(n2448) );
  NAND2X1 U4158 ( .A(\Mem[5][2] ), .B(n6613), .Y(n2167) );
  OAI21X1 U4159 ( .A(n6479), .B(n6609), .C(n2168), .Y(n2449) );
  NAND2X1 U4160 ( .A(\Mem[5][3] ), .B(n6612), .Y(n2168) );
  OAI21X1 U4161 ( .A(n6474), .B(n6609), .C(n2169), .Y(n2450) );
  NAND2X1 U4162 ( .A(\Mem[5][4] ), .B(n6613), .Y(n2169) );
  OAI21X1 U4163 ( .A(n6469), .B(n6609), .C(n2170), .Y(n2451) );
  NAND2X1 U4164 ( .A(\Mem[5][5] ), .B(n6612), .Y(n2170) );
  OAI21X1 U4165 ( .A(n6464), .B(n6609), .C(n2171), .Y(n2452) );
  NAND2X1 U4166 ( .A(\Mem[5][6] ), .B(n6612), .Y(n2171) );
  OAI21X1 U4167 ( .A(n6459), .B(n6609), .C(n2172), .Y(n2453) );
  NAND2X1 U4168 ( .A(\Mem[5][7] ), .B(n6612), .Y(n2172) );
  OAI21X1 U4169 ( .A(n6454), .B(n6609), .C(n2173), .Y(n2454) );
  NAND2X1 U4170 ( .A(\Mem[5][8] ), .B(n6612), .Y(n2173) );
  OAI21X1 U4171 ( .A(n6449), .B(n6609), .C(n2174), .Y(n2455) );
  NAND2X1 U4172 ( .A(\Mem[5][9] ), .B(n6612), .Y(n2174) );
  OAI21X1 U4173 ( .A(n6599), .B(n6609), .C(n2175), .Y(n2456) );
  NAND2X1 U4174 ( .A(\Mem[5][10] ), .B(n6612), .Y(n2175) );
  OAI21X1 U4175 ( .A(n6594), .B(n6609), .C(n2176), .Y(n2457) );
  NAND2X1 U4176 ( .A(\Mem[5][11] ), .B(n6612), .Y(n2176) );
  OAI21X1 U4177 ( .A(n6589), .B(n6609), .C(n2177), .Y(n2458) );
  NAND2X1 U4178 ( .A(\Mem[5][12] ), .B(n6612), .Y(n2177) );
  OAI21X1 U4179 ( .A(n6584), .B(n6610), .C(n2178), .Y(n2459) );
  NAND2X1 U4180 ( .A(\Mem[5][13] ), .B(n6612), .Y(n2178) );
  OAI21X1 U4181 ( .A(n6579), .B(n6610), .C(n2179), .Y(n2460) );
  NAND2X1 U4182 ( .A(\Mem[5][14] ), .B(n6612), .Y(n2179) );
  OAI21X1 U4183 ( .A(n6574), .B(n6610), .C(n2180), .Y(n2461) );
  NAND2X1 U4184 ( .A(\Mem[5][15] ), .B(n6611), .Y(n2180) );
  OAI21X1 U4185 ( .A(n6569), .B(n6610), .C(n2181), .Y(n2462) );
  NAND2X1 U4186 ( .A(\Mem[5][16] ), .B(n6612), .Y(n2181) );
  OAI21X1 U4187 ( .A(n6564), .B(n6610), .C(n2182), .Y(n2463) );
  NAND2X1 U4188 ( .A(\Mem[5][17] ), .B(n6611), .Y(n2182) );
  OAI21X1 U4189 ( .A(n6559), .B(n6610), .C(n2183), .Y(n2464) );
  NAND2X1 U4190 ( .A(\Mem[5][18] ), .B(n6611), .Y(n2183) );
  OAI21X1 U4191 ( .A(n6558), .B(n6610), .C(n2184), .Y(n2465) );
  NAND2X1 U4192 ( .A(\Mem[5][19] ), .B(n6611), .Y(n2184) );
  OAI21X1 U4194 ( .A(n6548), .B(n6610), .C(n2185), .Y(n2466) );
  NAND2X1 U4195 ( .A(\Mem[5][20] ), .B(n6611), .Y(n2185) );
  OAI21X1 U4197 ( .A(n6543), .B(n6610), .C(n2186), .Y(n2467) );
  NAND2X1 U4198 ( .A(\Mem[5][21] ), .B(n6611), .Y(n2186) );
  OAI21X1 U4200 ( .A(n6538), .B(n6610), .C(n2187), .Y(n2468) );
  NAND2X1 U4201 ( .A(\Mem[5][22] ), .B(n6612), .Y(n2187) );
  OAI21X1 U4203 ( .A(n6533), .B(n6611), .C(n2188), .Y(n2469) );
  NAND2X1 U4204 ( .A(\Mem[5][23] ), .B(n6611), .Y(n2188) );
  OAI21X1 U4206 ( .A(n6528), .B(n6610), .C(n2189), .Y(n2470) );
  NAND2X1 U4207 ( .A(\Mem[5][24] ), .B(n6612), .Y(n2189) );
  OAI21X1 U4209 ( .A(n6523), .B(n6611), .C(n2190), .Y(n2471) );
  NAND2X1 U4210 ( .A(\Mem[5][25] ), .B(n6612), .Y(n2190) );
  OAI21X1 U4212 ( .A(n6518), .B(n6611), .C(n2191), .Y(n2472) );
  NAND2X1 U4213 ( .A(\Mem[5][26] ), .B(n6612), .Y(n2191) );
  OAI21X1 U4215 ( .A(n6513), .B(n6611), .C(n2192), .Y(n2473) );
  NAND2X1 U4216 ( .A(\Mem[5][27] ), .B(n6612), .Y(n2192) );
  OAI21X1 U4218 ( .A(n6508), .B(n6611), .C(n2193), .Y(n2474) );
  NAND2X1 U4219 ( .A(\Mem[5][28] ), .B(n6612), .Y(n2193) );
  OAI21X1 U4221 ( .A(n6503), .B(n6611), .C(n2194), .Y(n2475) );
  NAND2X1 U4222 ( .A(\Mem[5][29] ), .B(n6612), .Y(n2194) );
  OAI21X1 U4224 ( .A(n6493), .B(n6611), .C(n2195), .Y(n2476) );
  NAND2X1 U4225 ( .A(\Mem[5][30] ), .B(n6613), .Y(n2195) );
  OAI21X1 U4227 ( .A(n6488), .B(n6611), .C(n2196), .Y(n2477) );
  NAND2X1 U4228 ( .A(\Mem[5][31] ), .B(n6613), .Y(n2196) );
  NAND2X1 U4229 ( .A(n7023), .B(n7004), .Y(n2164) );
  NAND3X1 U4231 ( .A(ADDR_WR[2]), .B(n7025), .C(ADDR_WR[0]), .Y(n2197) );
  OAI21X1 U4234 ( .A(n6924), .B(n6604), .C(n2198), .Y(n2478) );
  NAND2X1 U4235 ( .A(\Mem[6][0] ), .B(n6927), .Y(n2198) );
  OAI21X1 U4237 ( .A(n6925), .B(n6549), .C(n2199), .Y(n2479) );
  NAND2X1 U4238 ( .A(\Mem[6][1] ), .B(n6926), .Y(n2199) );
  OAI21X1 U4240 ( .A(n6925), .B(n6494), .C(n2200), .Y(n2480) );
  NAND2X1 U4241 ( .A(\Mem[6][2] ), .B(n6926), .Y(n2200) );
  OAI21X1 U4243 ( .A(n6925), .B(n6479), .C(n2201), .Y(n2481) );
  NAND2X1 U4244 ( .A(\Mem[6][3] ), .B(n6927), .Y(n2201) );
  OAI21X1 U4246 ( .A(n6925), .B(n6474), .C(n2202), .Y(n2482) );
  NAND2X1 U4247 ( .A(\Mem[6][4] ), .B(n6926), .Y(n2202) );
  OAI21X1 U4249 ( .A(n6925), .B(n6469), .C(n2203), .Y(n2483) );
  NAND2X1 U4250 ( .A(\Mem[6][5] ), .B(n6926), .Y(n2203) );
  OAI21X1 U4252 ( .A(n6925), .B(n6464), .C(n2204), .Y(n2484) );
  NAND2X1 U4253 ( .A(\Mem[6][6] ), .B(n6926), .Y(n2204) );
  OAI21X1 U4255 ( .A(n6925), .B(n6459), .C(n2205), .Y(n2485) );
  NAND2X1 U4256 ( .A(\Mem[6][7] ), .B(n6926), .Y(n2205) );
  OAI21X1 U4258 ( .A(n6925), .B(n6454), .C(n2206), .Y(n2486) );
  NAND2X1 U4259 ( .A(\Mem[6][8] ), .B(n6926), .Y(n2206) );
  OAI21X1 U4261 ( .A(n6925), .B(n6449), .C(n2207), .Y(n2487) );
  NAND2X1 U4262 ( .A(\Mem[6][9] ), .B(n6927), .Y(n2207) );
  OAI21X1 U4264 ( .A(n6925), .B(n6599), .C(n2208), .Y(n2488) );
  NAND2X1 U4265 ( .A(\Mem[6][10] ), .B(n6926), .Y(n2208) );
  OAI21X1 U4267 ( .A(n6925), .B(n6594), .C(n2209), .Y(n2489) );
  NAND2X1 U4268 ( .A(\Mem[6][11] ), .B(n6926), .Y(n2209) );
  OAI21X1 U4270 ( .A(n6926), .B(n6589), .C(n2210), .Y(n2490) );
  NAND2X1 U4271 ( .A(\Mem[6][12] ), .B(n6927), .Y(n2210) );
  OAI21X1 U4273 ( .A(n6926), .B(n6584), .C(n2211), .Y(n2491) );
  NAND2X1 U4274 ( .A(\Mem[6][13] ), .B(n6927), .Y(n2211) );
  OAI21X1 U4276 ( .A(n6925), .B(n6579), .C(n2212), .Y(n2492) );
  NAND2X1 U4277 ( .A(\Mem[6][14] ), .B(n6927), .Y(n2212) );
  OAI21X1 U4279 ( .A(n6926), .B(n6574), .C(n2213), .Y(n2493) );
  NAND2X1 U4280 ( .A(\Mem[6][15] ), .B(n6927), .Y(n2213) );
  OAI21X1 U4282 ( .A(n6926), .B(n6569), .C(n2214), .Y(n2494) );
  NAND2X1 U4283 ( .A(\Mem[6][16] ), .B(n6927), .Y(n2214) );
  OAI21X1 U4285 ( .A(n6926), .B(n6564), .C(n2215), .Y(n2495) );
  NAND2X1 U4286 ( .A(\Mem[6][17] ), .B(n6928), .Y(n2215) );
  OAI21X1 U4288 ( .A(n6926), .B(n6559), .C(n2216), .Y(n2496) );
  NAND2X1 U4289 ( .A(\Mem[6][18] ), .B(n6928), .Y(n2216) );
  NAND2X1 U4291 ( .A(n7024), .B(n7004), .Y(n1) );
  NAND3X1 U4293 ( .A(n7015), .B(n7014), .C(n81), .Y(n2217) );
  NOR2X1 U4294 ( .A(n1957), .B(ADDR_WR[5]), .Y(n355) );
  NAND3X1 U4295 ( .A(WR), .B(n7012), .C(n2219), .Y(n1957) );
  NOR2X1 U4296 ( .A(ADDR_WR[8]), .B(ADDR_WR[7]), .Y(n2219) );
  NAND3X1 U4301 ( .A(ADDR_WR[1]), .B(n7026), .C(ADDR_WR[2]), .Y(n2220) );
  DFFSR \DOUT_reg[1]  ( .D(n6970), .CLK(clk), .R(n7027), .S(1'b1), .Q(DOUT[1])
         );
  DFFSR \DOUT_reg[5]  ( .D(n6966), .CLK(clk), .R(n7027), .S(1'b1), .Q(DOUT[5])
         );
  DFFSR \DOUT_reg[4]  ( .D(n6967), .CLK(clk), .R(n7027), .S(1'b1), .Q(DOUT[4])
         );
  DFFSR \DOUT_reg[3]  ( .D(n6968), .CLK(clk), .R(n7027), .S(1'b1), .Q(DOUT[3])
         );
  DFFSR \DOUT_reg[2]  ( .D(n6969), .CLK(clk), .R(n7027), .S(1'b1), .Q(DOUT[2])
         );
  DFFSR \DOUT_reg[18]  ( .D(n6953), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[18]) );
  DFFSR \DOUT_reg[17]  ( .D(n6954), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[17]) );
  DFFSR \DOUT_reg[16]  ( .D(n6955), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[16]) );
  DFFSR \DOUT_reg[15]  ( .D(n6956), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[15]) );
  DFFSR \DOUT_reg[14]  ( .D(n6957), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[14]) );
  DFFSR \DOUT_reg[13]  ( .D(n6958), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[13]) );
  DFFSR \DOUT_reg[12]  ( .D(n6959), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[12]) );
  DFFSR \DOUT_reg[11]  ( .D(n6960), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[11]) );
  DFFSR \DOUT_reg[10]  ( .D(n6961), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[10]) );
  DFFSR \DOUT_reg[9]  ( .D(n6962), .CLK(clk), .R(n7027), .S(1'b1), .Q(DOUT[9])
         );
  DFFSR \DOUT_reg[8]  ( .D(n6963), .CLK(clk), .R(n7027), .S(1'b1), .Q(DOUT[8])
         );
  DFFSR \DOUT_reg[7]  ( .D(n6964), .CLK(clk), .R(n7027), .S(1'b1), .Q(DOUT[7])
         );
  DFFSR \DOUT_reg[6]  ( .D(n6965), .CLK(clk), .R(n7027), .S(1'b1), .Q(DOUT[6])
         );
  DFFSR \DOUT_reg[31]  ( .D(n6940), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[31]) );
  DFFSR \DOUT_reg[30]  ( .D(n6941), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[30]) );
  DFFSR \DOUT_reg[29]  ( .D(n6942), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[29]) );
  DFFSR \DOUT_reg[28]  ( .D(n6943), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[28]) );
  DFFSR \DOUT_reg[27]  ( .D(n6944), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[27]) );
  DFFSR \DOUT_reg[26]  ( .D(n6945), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[26]) );
  DFFSR \DOUT_reg[25]  ( .D(n6946), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[25]) );
  DFFSR \DOUT_reg[24]  ( .D(n6947), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[24]) );
  DFFSR \DOUT_reg[23]  ( .D(n6948), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[23]) );
  DFFSR \DOUT_reg[22]  ( .D(n6949), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[22]) );
  DFFSR \DOUT_reg[21]  ( .D(n6950), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[21]) );
  DFFSR \DOUT_reg[20]  ( .D(n6951), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[20]) );
  DFFSR \DOUT_reg[19]  ( .D(n6952), .CLK(clk), .R(n7027), .S(1'b1), .Q(
        DOUT[19]) );
  DFFSR \DOUT_reg[0]  ( .D(n6971), .CLK(clk), .R(n7027), .S(1'b1), .Q(DOUT[0])
         );
  INVX4 U613 ( .A(reset), .Y(n7027) );
  BUFX2 U3799 ( .A(n1156), .Y(n80) );
  NOR2X1 U3801 ( .A(n1957), .B(ADDR_WR[5]), .Y(n81) );
  BUFX2 U3803 ( .A(n6360), .Y(n6362) );
  BUFX2 U3805 ( .A(n6359), .Y(n6365) );
  BUFX2 U3807 ( .A(n6359), .Y(n6364) );
  BUFX2 U3809 ( .A(n6360), .Y(n6363) );
  BUFX2 U3811 ( .A(n6358), .Y(n6367) );
  BUFX2 U3813 ( .A(n6359), .Y(n6366) );
  BUFX2 U3814 ( .A(n6357), .Y(n6370) );
  BUFX2 U3816 ( .A(n6358), .Y(n6369) );
  BUFX2 U3882 ( .A(n6358), .Y(n6368) );
  BUFX2 U3949 ( .A(n6357), .Y(n6372) );
  BUFX2 U4016 ( .A(n6357), .Y(n6371) );
  BUFX2 U4083 ( .A(n6356), .Y(n6375) );
  BUFX2 U4085 ( .A(n6356), .Y(n6374) );
  BUFX2 U4151 ( .A(n6356), .Y(n6373) );
  BUFX2 U4193 ( .A(n6355), .Y(n6377) );
  BUFX2 U4196 ( .A(n6355), .Y(n6376) );
  BUFX2 U4199 ( .A(n6354), .Y(n6379) );
  BUFX2 U4202 ( .A(n6355), .Y(n6378) );
  BUFX2 U4205 ( .A(n6353), .Y(n6382) );
  BUFX2 U4208 ( .A(n6354), .Y(n6381) );
  BUFX2 U4211 ( .A(n6354), .Y(n6380) );
  BUFX2 U4214 ( .A(n6353), .Y(n6384) );
  BUFX2 U4217 ( .A(n6353), .Y(n6383) );
  BUFX2 U4220 ( .A(n6352), .Y(n6387) );
  BUFX2 U4223 ( .A(n6352), .Y(n6386) );
  BUFX2 U4226 ( .A(n6352), .Y(n6385) );
  BUFX2 U4230 ( .A(n6351), .Y(n6389) );
  BUFX2 U4232 ( .A(n6351), .Y(n6388) );
  BUFX2 U4233 ( .A(n6350), .Y(n6392) );
  BUFX2 U4236 ( .A(n6350), .Y(n6391) );
  BUFX2 U4239 ( .A(n6351), .Y(n6390) );
  BUFX2 U4242 ( .A(n6349), .Y(n6394) );
  BUFX2 U4245 ( .A(n6350), .Y(n6393) );
  BUFX2 U4248 ( .A(n6348), .Y(n6397) );
  BUFX2 U4251 ( .A(n6349), .Y(n6396) );
  BUFX2 U4254 ( .A(n6349), .Y(n6395) );
  BUFX2 U4257 ( .A(n6348), .Y(n6399) );
  BUFX2 U4260 ( .A(n6348), .Y(n6398) );
  BUFX2 U4263 ( .A(n6347), .Y(n6402) );
  BUFX2 U4266 ( .A(n6347), .Y(n6401) );
  BUFX2 U4269 ( .A(n6347), .Y(n6400) );
  BUFX2 U4272 ( .A(n6346), .Y(n6404) );
  BUFX2 U4275 ( .A(n6346), .Y(n6403) );
  BUFX2 U4278 ( .A(n6345), .Y(n6407) );
  BUFX2 U4281 ( .A(n6345), .Y(n6406) );
  BUFX2 U4284 ( .A(n6346), .Y(n6405) );
  BUFX2 U4287 ( .A(n6344), .Y(n6409) );
  BUFX2 U4290 ( .A(n6345), .Y(n6408) );
  BUFX2 U4292 ( .A(n6344), .Y(n6411) );
  BUFX2 U4297 ( .A(n6344), .Y(n6410) );
  BUFX2 U4298 ( .A(n6343), .Y(n6414) );
  BUFX2 U4299 ( .A(n6343), .Y(n6413) );
  BUFX2 U4300 ( .A(n6343), .Y(n6412) );
  BUFX2 U4302 ( .A(n6342), .Y(n6416) );
  BUFX2 U4303 ( .A(n6342), .Y(n6415) );
  BUFX2 U4304 ( .A(n6341), .Y(n6419) );
  BUFX2 U4305 ( .A(n6341), .Y(n6418) );
  BUFX2 U4306 ( .A(n6342), .Y(n6417) );
  BUFX2 U4307 ( .A(n6340), .Y(n6421) );
  BUFX2 U4308 ( .A(n6341), .Y(n6420) );
  BUFX2 U4309 ( .A(n6339), .Y(n6424) );
  BUFX2 U4310 ( .A(n6340), .Y(n6423) );
  BUFX2 U4311 ( .A(n6340), .Y(n6422) );
  BUFX2 U4312 ( .A(n6339), .Y(n6426) );
  BUFX2 U4313 ( .A(n6339), .Y(n6425) );
  BUFX2 U4314 ( .A(n6338), .Y(n6429) );
  BUFX2 U4315 ( .A(n6338), .Y(n6428) );
  BUFX2 U4316 ( .A(n6338), .Y(n6427) );
  BUFX2 U4317 ( .A(n6337), .Y(n6431) );
  BUFX2 U4318 ( .A(n6337), .Y(n6430) );
  BUFX2 U4319 ( .A(n6336), .Y(n6434) );
  BUFX2 U4320 ( .A(n6336), .Y(n6433) );
  BUFX2 U4321 ( .A(n6337), .Y(n6432) );
  BUFX2 U4322 ( .A(n6335), .Y(n6436) );
  BUFX2 U4323 ( .A(n6336), .Y(n6435) );
  BUFX2 U4324 ( .A(n6335), .Y(n6438) );
  BUFX2 U4325 ( .A(n6335), .Y(n6437) );
  BUFX2 U4326 ( .A(n6288), .Y(n6291) );
  BUFX2 U4327 ( .A(n6288), .Y(n6290) );
  BUFX2 U4328 ( .A(n6287), .Y(n6292) );
  BUFX2 U4329 ( .A(n6287), .Y(n6293) );
  BUFX2 U4330 ( .A(n6287), .Y(n6294) );
  BUFX2 U4331 ( .A(n6286), .Y(n6296) );
  BUFX2 U4332 ( .A(n6286), .Y(n6295) );
  BUFX2 U4333 ( .A(n6286), .Y(n6297) );
  BUFX2 U4334 ( .A(n6285), .Y(n6298) );
  BUFX2 U4335 ( .A(n6285), .Y(n6299) );
  BUFX2 U4336 ( .A(n6285), .Y(n6300) );
  BUFX2 U4337 ( .A(n6284), .Y(n6302) );
  BUFX2 U4338 ( .A(n6284), .Y(n6301) );
  BUFX2 U4339 ( .A(n6284), .Y(n6303) );
  BUFX2 U4340 ( .A(n6283), .Y(n6304) );
  BUFX2 U4341 ( .A(n6283), .Y(n6305) );
  BUFX2 U4342 ( .A(n6282), .Y(n6307) );
  BUFX2 U4343 ( .A(n6283), .Y(n6306) );
  BUFX2 U4344 ( .A(n6282), .Y(n6308) );
  BUFX2 U4345 ( .A(n6282), .Y(n6309) );
  BUFX2 U4346 ( .A(n6281), .Y(n6310) );
  BUFX2 U4347 ( .A(n6281), .Y(n6312) );
  BUFX2 U4348 ( .A(n6281), .Y(n6311) );
  BUFX2 U4349 ( .A(n6280), .Y(n6313) );
  BUFX2 U4350 ( .A(n6280), .Y(n6314) );
  BUFX2 U4351 ( .A(n6280), .Y(n6315) );
  BUFX2 U4352 ( .A(n6279), .Y(n6316) );
  BUFX2 U4353 ( .A(n6279), .Y(n6318) );
  BUFX2 U4354 ( .A(n6279), .Y(n6317) );
  BUFX2 U4355 ( .A(n6278), .Y(n6319) );
  BUFX2 U4356 ( .A(n6278), .Y(n6320) );
  BUFX2 U4357 ( .A(n6278), .Y(n6321) );
  BUFX2 U4358 ( .A(n6277), .Y(n6323) );
  BUFX2 U4359 ( .A(n6277), .Y(n6322) );
  BUFX2 U4360 ( .A(n6277), .Y(n6324) );
  BUFX2 U4361 ( .A(n6276), .Y(n6325) );
  BUFX2 U4362 ( .A(n6276), .Y(n6326) );
  BUFX2 U4363 ( .A(n6276), .Y(n6327) );
  BUFX2 U4364 ( .A(n6360), .Y(n6361) );
  INVX2 U4365 ( .A(n6934), .Y(n6929) );
  INVX2 U4366 ( .A(n6933), .Y(n6930) );
  BUFX2 U4367 ( .A(n6288), .Y(n6289) );
  INVX2 U4368 ( .A(n6932), .Y(n6931) );
  BUFX2 U4369 ( .A(n1991), .Y(n6636) );
  BUFX2 U4370 ( .A(n890), .Y(n6796) );
  BUFX2 U4371 ( .A(n1991), .Y(n6637) );
  BUFX2 U4372 ( .A(n890), .Y(n6797) );
  BUFX2 U4373 ( .A(n1991), .Y(n6634) );
  BUFX2 U4374 ( .A(n1991), .Y(n6635) );
  BUFX2 U4375 ( .A(n890), .Y(n6794) );
  BUFX2 U4376 ( .A(n890), .Y(n6795) );
  BUFX2 U4377 ( .A(n1991), .Y(n6638) );
  BUFX2 U4378 ( .A(n890), .Y(n6798) );
  BUFX2 U4379 ( .A(n6269), .Y(n6250) );
  BUFX2 U4380 ( .A(n6269), .Y(n6251) );
  BUFX2 U4381 ( .A(n6269), .Y(n6252) );
  BUFX2 U4382 ( .A(n6270), .Y(n6253) );
  BUFX2 U4383 ( .A(n6270), .Y(n6254) );
  BUFX2 U4384 ( .A(n6270), .Y(n6255) );
  BUFX2 U4385 ( .A(n6271), .Y(n6256) );
  BUFX2 U4386 ( .A(n6271), .Y(n6257) );
  BUFX2 U4387 ( .A(n6271), .Y(n6258) );
  BUFX2 U4388 ( .A(n6272), .Y(n6259) );
  BUFX2 U4389 ( .A(n6272), .Y(n6260) );
  BUFX2 U4390 ( .A(n6272), .Y(n6261) );
  BUFX2 U4391 ( .A(n6273), .Y(n6262) );
  BUFX2 U4392 ( .A(n6273), .Y(n6263) );
  BUFX2 U4393 ( .A(n6273), .Y(n6264) );
  BUFX2 U4394 ( .A(n6274), .Y(n6265) );
  BUFX2 U4395 ( .A(n6274), .Y(n6266) );
  BUFX2 U4396 ( .A(n6274), .Y(n6267) );
  BUFX2 U4397 ( .A(n6268), .Y(n6249) );
  BUFX2 U4398 ( .A(n6334), .Y(n6439) );
  BUFX2 U4399 ( .A(n6440), .Y(n6334) );
  BUFX2 U4400 ( .A(n6275), .Y(n6328) );
  BUFX2 U4401 ( .A(n6329), .Y(n6275) );
  BUFX2 U4402 ( .A(n6268), .Y(n6248) );
  BUFX2 U4403 ( .A(n6939), .Y(n6934) );
  BUFX2 U4404 ( .A(n6938), .Y(n6933) );
  BUFX2 U4405 ( .A(n6939), .Y(n6932) );
  BUFX2 U4406 ( .A(n6939), .Y(n6937) );
  BUFX2 U4407 ( .A(n6939), .Y(n6936) );
  BUFX2 U4408 ( .A(n6939), .Y(n6935) );
  BUFX2 U4409 ( .A(n6329), .Y(n6276) );
  BUFX2 U4410 ( .A(n6448), .Y(n6360) );
  BUFX2 U4411 ( .A(n6448), .Y(n6359) );
  BUFX2 U4412 ( .A(n6448), .Y(n6358) );
  BUFX2 U4413 ( .A(n6447), .Y(n6357) );
  BUFX2 U4414 ( .A(n6447), .Y(n6356) );
  BUFX2 U4415 ( .A(n6447), .Y(n6355) );
  BUFX2 U4416 ( .A(n6446), .Y(n6354) );
  BUFX2 U4417 ( .A(n6446), .Y(n6353) );
  BUFX2 U4418 ( .A(n6446), .Y(n6352) );
  BUFX2 U4419 ( .A(n6445), .Y(n6351) );
  BUFX2 U4420 ( .A(n6445), .Y(n6350) );
  BUFX2 U4421 ( .A(n6445), .Y(n6349) );
  BUFX2 U4422 ( .A(n6444), .Y(n6348) );
  BUFX2 U4423 ( .A(n6444), .Y(n6347) );
  BUFX2 U4424 ( .A(n6444), .Y(n6346) );
  BUFX2 U4425 ( .A(n6443), .Y(n6345) );
  BUFX2 U4426 ( .A(n6443), .Y(n6344) );
  BUFX2 U4427 ( .A(n6443), .Y(n6343) );
  BUFX2 U4428 ( .A(n6442), .Y(n6342) );
  BUFX2 U4429 ( .A(n6442), .Y(n6341) );
  BUFX2 U4430 ( .A(n6442), .Y(n6340) );
  BUFX2 U4431 ( .A(n6441), .Y(n6339) );
  BUFX2 U4432 ( .A(n6441), .Y(n6338) );
  BUFX2 U4433 ( .A(n6441), .Y(n6337) );
  BUFX2 U4434 ( .A(n6440), .Y(n6336) );
  BUFX2 U4435 ( .A(n6440), .Y(n6335) );
  BUFX2 U4436 ( .A(n6333), .Y(n6288) );
  BUFX2 U4437 ( .A(n6333), .Y(n6287) );
  BUFX2 U4438 ( .A(n6333), .Y(n6286) );
  BUFX2 U4439 ( .A(n6332), .Y(n6285) );
  BUFX2 U4440 ( .A(n6332), .Y(n6284) );
  BUFX2 U4441 ( .A(n6332), .Y(n6283) );
  BUFX2 U4442 ( .A(n6331), .Y(n6282) );
  BUFX2 U4443 ( .A(n6331), .Y(n6281) );
  BUFX2 U4444 ( .A(n6331), .Y(n6280) );
  BUFX2 U4445 ( .A(n6330), .Y(n6279) );
  BUFX2 U4446 ( .A(n6330), .Y(n6278) );
  BUFX2 U4447 ( .A(n6330), .Y(n6277) );
  BUFX2 U4448 ( .A(n6939), .Y(n6938) );
  BUFX2 U4449 ( .A(n28), .Y(n6920) );
  BUFX2 U4450 ( .A(n1), .Y(n6925) );
  BUFX2 U4451 ( .A(n1), .Y(n6924) );
  BUFX2 U4452 ( .A(n2096), .Y(n6621) );
  BUFX2 U4453 ( .A(n2164), .Y(n6611) );
  BUFX2 U4454 ( .A(n185), .Y(n6901) );
  BUFX2 U4455 ( .A(n253), .Y(n6891) );
  BUFX2 U4456 ( .A(n287), .Y(n6886) );
  BUFX2 U4457 ( .A(n321), .Y(n6881) );
  BUFX2 U4458 ( .A(n624), .Y(n6836) );
  BUFX2 U4459 ( .A(n658), .Y(n6831) );
  BUFX2 U4460 ( .A(n691), .Y(n6826) );
  BUFX2 U4461 ( .A(n724), .Y(n6821) );
  BUFX2 U4462 ( .A(n757), .Y(n6816) );
  BUFX2 U4463 ( .A(n790), .Y(n6811) );
  BUFX2 U4464 ( .A(n823), .Y(n6806) );
  BUFX2 U4465 ( .A(n856), .Y(n6801) );
  BUFX2 U4466 ( .A(n1157), .Y(n6756) );
  BUFX2 U4467 ( .A(n1191), .Y(n6751) );
  BUFX2 U4468 ( .A(n1224), .Y(n6746) );
  BUFX2 U4469 ( .A(n1257), .Y(n6741) );
  BUFX2 U4470 ( .A(n1290), .Y(n6736) );
  BUFX2 U4471 ( .A(n1323), .Y(n6731) );
  BUFX2 U4472 ( .A(n1356), .Y(n6726) );
  BUFX2 U4473 ( .A(n1389), .Y(n6721) );
  BUFX2 U4474 ( .A(n1423), .Y(n6716) );
  BUFX2 U4475 ( .A(n1457), .Y(n6711) );
  BUFX2 U4476 ( .A(n1490), .Y(n6706) );
  BUFX2 U4477 ( .A(n1523), .Y(n6701) );
  BUFX2 U4478 ( .A(n1556), .Y(n6696) );
  BUFX2 U4479 ( .A(n1589), .Y(n6691) );
  BUFX2 U4480 ( .A(n1622), .Y(n6686) );
  BUFX2 U4481 ( .A(n1655), .Y(n6681) );
  BUFX2 U4482 ( .A(n1689), .Y(n6676) );
  BUFX2 U4483 ( .A(n1723), .Y(n6671) );
  BUFX2 U4484 ( .A(n1756), .Y(n6666) );
  BUFX2 U4485 ( .A(n1789), .Y(n6661) );
  BUFX2 U4486 ( .A(n1822), .Y(n6656) );
  BUFX2 U4487 ( .A(n1855), .Y(n6651) );
  BUFX2 U4488 ( .A(n1888), .Y(n6646) );
  BUFX2 U4489 ( .A(n1921), .Y(n6641) );
  BUFX2 U4490 ( .A(n2028), .Y(n6631) );
  BUFX2 U4491 ( .A(n2062), .Y(n6626) );
  BUFX2 U4492 ( .A(n2130), .Y(n6616) );
  BUFX2 U4493 ( .A(n82), .Y(n6916) );
  BUFX2 U4494 ( .A(n117), .Y(n6911) );
  BUFX2 U4495 ( .A(n151), .Y(n6906) );
  BUFX2 U4496 ( .A(n219), .Y(n6896) );
  BUFX2 U4497 ( .A(n357), .Y(n6876) );
  BUFX2 U4498 ( .A(n391), .Y(n6871) );
  BUFX2 U4499 ( .A(n424), .Y(n6866) );
  BUFX2 U4500 ( .A(n457), .Y(n6861) );
  BUFX2 U4501 ( .A(n490), .Y(n6856) );
  BUFX2 U4502 ( .A(n523), .Y(n6851) );
  BUFX2 U4503 ( .A(n556), .Y(n6846) );
  BUFX2 U4504 ( .A(n589), .Y(n6841) );
  BUFX2 U4505 ( .A(n924), .Y(n6791) );
  BUFX2 U4506 ( .A(n957), .Y(n6786) );
  BUFX2 U4507 ( .A(n990), .Y(n6781) );
  BUFX2 U4508 ( .A(n1023), .Y(n6776) );
  BUFX2 U4509 ( .A(n1056), .Y(n6771) );
  BUFX2 U4510 ( .A(n1089), .Y(n6766) );
  BUFX2 U4511 ( .A(n1122), .Y(n6761) );
  BUFX2 U4512 ( .A(n2096), .Y(n6622) );
  BUFX2 U4513 ( .A(n2164), .Y(n6612) );
  BUFX2 U4514 ( .A(n28), .Y(n6922) );
  BUFX2 U4515 ( .A(n185), .Y(n6902) );
  BUFX2 U4516 ( .A(n253), .Y(n6892) );
  BUFX2 U4517 ( .A(n287), .Y(n6887) );
  BUFX2 U4518 ( .A(n321), .Y(n6882) );
  BUFX2 U4519 ( .A(n1224), .Y(n6747) );
  BUFX2 U4520 ( .A(n1257), .Y(n6742) );
  BUFX2 U4521 ( .A(n1290), .Y(n6737) );
  BUFX2 U4522 ( .A(n1323), .Y(n6732) );
  BUFX2 U4523 ( .A(n1356), .Y(n6727) );
  BUFX2 U4524 ( .A(n1389), .Y(n6722) );
  BUFX2 U4525 ( .A(n1423), .Y(n6717) );
  BUFX2 U4526 ( .A(n1457), .Y(n6712) );
  BUFX2 U4527 ( .A(n1490), .Y(n6707) );
  BUFX2 U4528 ( .A(n1523), .Y(n6702) );
  BUFX2 U4529 ( .A(n1556), .Y(n6697) );
  BUFX2 U4530 ( .A(n1589), .Y(n6692) );
  BUFX2 U4531 ( .A(n1622), .Y(n6687) );
  BUFX2 U4532 ( .A(n1655), .Y(n6682) );
  BUFX2 U4533 ( .A(n1689), .Y(n6677) );
  BUFX2 U4534 ( .A(n1723), .Y(n6672) );
  BUFX2 U4535 ( .A(n1756), .Y(n6667) );
  BUFX2 U4536 ( .A(n1789), .Y(n6662) );
  BUFX2 U4537 ( .A(n1822), .Y(n6657) );
  BUFX2 U4538 ( .A(n1855), .Y(n6652) );
  BUFX2 U4539 ( .A(n1888), .Y(n6647) );
  BUFX2 U4540 ( .A(n1921), .Y(n6642) );
  BUFX2 U4541 ( .A(n2028), .Y(n6632) );
  BUFX2 U4542 ( .A(n2062), .Y(n6627) );
  BUFX2 U4543 ( .A(n2130), .Y(n6617) );
  BUFX2 U4544 ( .A(n82), .Y(n6917) );
  BUFX2 U4545 ( .A(n117), .Y(n6912) );
  BUFX2 U4546 ( .A(n151), .Y(n6907) );
  BUFX2 U4547 ( .A(n219), .Y(n6897) );
  BUFX2 U4548 ( .A(n357), .Y(n6877) );
  BUFX2 U4549 ( .A(n391), .Y(n6872) );
  BUFX2 U4550 ( .A(n424), .Y(n6867) );
  BUFX2 U4551 ( .A(n457), .Y(n6862) );
  BUFX2 U4552 ( .A(n490), .Y(n6857) );
  BUFX2 U4553 ( .A(n523), .Y(n6852) );
  BUFX2 U4554 ( .A(n556), .Y(n6847) );
  BUFX2 U4555 ( .A(n589), .Y(n6842) );
  BUFX2 U4556 ( .A(n624), .Y(n6837) );
  BUFX2 U4557 ( .A(n658), .Y(n6832) );
  BUFX2 U4558 ( .A(n691), .Y(n6827) );
  BUFX2 U4559 ( .A(n724), .Y(n6822) );
  BUFX2 U4560 ( .A(n757), .Y(n6817) );
  BUFX2 U4561 ( .A(n790), .Y(n6812) );
  BUFX2 U4562 ( .A(n823), .Y(n6807) );
  BUFX2 U4563 ( .A(n856), .Y(n6802) );
  BUFX2 U4564 ( .A(n1157), .Y(n6757) );
  BUFX2 U4565 ( .A(n1191), .Y(n6752) );
  BUFX2 U4566 ( .A(n924), .Y(n6792) );
  BUFX2 U4567 ( .A(n957), .Y(n6787) );
  BUFX2 U4568 ( .A(n990), .Y(n6782) );
  BUFX2 U4569 ( .A(n1023), .Y(n6777) );
  BUFX2 U4570 ( .A(n1056), .Y(n6772) );
  BUFX2 U4571 ( .A(n1089), .Y(n6767) );
  BUFX2 U4572 ( .A(n1122), .Y(n6762) );
  BUFX2 U4573 ( .A(n28), .Y(n6921) );
  BUFX2 U4574 ( .A(n2096), .Y(n6619) );
  BUFX2 U4575 ( .A(n2096), .Y(n6620) );
  BUFX2 U4576 ( .A(n2164), .Y(n6609) );
  BUFX2 U4577 ( .A(n2164), .Y(n6610) );
  BUFX2 U4578 ( .A(n28), .Y(n6919) );
  BUFX2 U4579 ( .A(n185), .Y(n6899) );
  BUFX2 U4580 ( .A(n185), .Y(n6900) );
  BUFX2 U4581 ( .A(n253), .Y(n6889) );
  BUFX2 U4582 ( .A(n253), .Y(n6890) );
  BUFX2 U4583 ( .A(n287), .Y(n6884) );
  BUFX2 U4584 ( .A(n287), .Y(n6885) );
  BUFX2 U4585 ( .A(n321), .Y(n6879) );
  BUFX2 U4586 ( .A(n321), .Y(n6880) );
  BUFX2 U4587 ( .A(n624), .Y(n6834) );
  BUFX2 U4588 ( .A(n624), .Y(n6835) );
  BUFX2 U4589 ( .A(n658), .Y(n6829) );
  BUFX2 U4590 ( .A(n658), .Y(n6830) );
  BUFX2 U4591 ( .A(n691), .Y(n6824) );
  BUFX2 U4592 ( .A(n691), .Y(n6825) );
  BUFX2 U4593 ( .A(n724), .Y(n6819) );
  BUFX2 U4594 ( .A(n724), .Y(n6820) );
  BUFX2 U4595 ( .A(n757), .Y(n6814) );
  BUFX2 U4596 ( .A(n757), .Y(n6815) );
  BUFX2 U4597 ( .A(n790), .Y(n6809) );
  BUFX2 U4598 ( .A(n790), .Y(n6810) );
  BUFX2 U4599 ( .A(n823), .Y(n6804) );
  BUFX2 U4600 ( .A(n823), .Y(n6805) );
  BUFX2 U4601 ( .A(n856), .Y(n6799) );
  BUFX2 U4602 ( .A(n856), .Y(n6800) );
  BUFX2 U4603 ( .A(n1157), .Y(n6754) );
  BUFX2 U4604 ( .A(n1157), .Y(n6755) );
  BUFX2 U4605 ( .A(n1191), .Y(n6749) );
  BUFX2 U4606 ( .A(n1191), .Y(n6750) );
  BUFX2 U4607 ( .A(n1224), .Y(n6744) );
  BUFX2 U4608 ( .A(n1224), .Y(n6745) );
  BUFX2 U4609 ( .A(n1257), .Y(n6739) );
  BUFX2 U4610 ( .A(n1257), .Y(n6740) );
  BUFX2 U4611 ( .A(n1290), .Y(n6734) );
  BUFX2 U4612 ( .A(n1290), .Y(n6735) );
  BUFX2 U4613 ( .A(n1323), .Y(n6729) );
  BUFX2 U4614 ( .A(n1323), .Y(n6730) );
  BUFX2 U4615 ( .A(n1356), .Y(n6724) );
  BUFX2 U4616 ( .A(n1356), .Y(n6725) );
  BUFX2 U4617 ( .A(n1389), .Y(n6719) );
  BUFX2 U4618 ( .A(n1389), .Y(n6720) );
  BUFX2 U4619 ( .A(n1423), .Y(n6714) );
  BUFX2 U4620 ( .A(n1423), .Y(n6715) );
  BUFX2 U4621 ( .A(n1457), .Y(n6709) );
  BUFX2 U4622 ( .A(n1457), .Y(n6710) );
  BUFX2 U4623 ( .A(n1490), .Y(n6704) );
  BUFX2 U4624 ( .A(n1490), .Y(n6705) );
  BUFX2 U4625 ( .A(n1523), .Y(n6699) );
  BUFX2 U4626 ( .A(n1523), .Y(n6700) );
  BUFX2 U4627 ( .A(n1556), .Y(n6694) );
  BUFX2 U4628 ( .A(n1556), .Y(n6695) );
  BUFX2 U4629 ( .A(n1589), .Y(n6689) );
  BUFX2 U4630 ( .A(n1589), .Y(n6690) );
  BUFX2 U4631 ( .A(n1622), .Y(n6684) );
  BUFX2 U4632 ( .A(n1622), .Y(n6685) );
  BUFX2 U4633 ( .A(n1655), .Y(n6679) );
  BUFX2 U4634 ( .A(n1655), .Y(n6680) );
  BUFX2 U4635 ( .A(n1689), .Y(n6674) );
  BUFX2 U4636 ( .A(n1689), .Y(n6675) );
  BUFX2 U4637 ( .A(n1723), .Y(n6669) );
  BUFX2 U4638 ( .A(n1723), .Y(n6670) );
  BUFX2 U4639 ( .A(n1756), .Y(n6664) );
  BUFX2 U4640 ( .A(n1756), .Y(n6665) );
  BUFX2 U4641 ( .A(n1789), .Y(n6659) );
  BUFX2 U4642 ( .A(n1789), .Y(n6660) );
  BUFX2 U4643 ( .A(n1822), .Y(n6654) );
  BUFX2 U4644 ( .A(n1822), .Y(n6655) );
  BUFX2 U4645 ( .A(n1855), .Y(n6649) );
  BUFX2 U4646 ( .A(n1855), .Y(n6650) );
  BUFX2 U4647 ( .A(n1888), .Y(n6644) );
  BUFX2 U4648 ( .A(n1888), .Y(n6645) );
  BUFX2 U4649 ( .A(n1921), .Y(n6639) );
  BUFX2 U4650 ( .A(n1921), .Y(n6640) );
  BUFX2 U4651 ( .A(n2028), .Y(n6629) );
  BUFX2 U4652 ( .A(n2028), .Y(n6630) );
  BUFX2 U4653 ( .A(n2062), .Y(n6624) );
  BUFX2 U4654 ( .A(n2062), .Y(n6625) );
  BUFX2 U4655 ( .A(n2130), .Y(n6614) );
  BUFX2 U4656 ( .A(n2130), .Y(n6615) );
  BUFX2 U4657 ( .A(n82), .Y(n6914) );
  BUFX2 U4658 ( .A(n82), .Y(n6915) );
  BUFX2 U4659 ( .A(n117), .Y(n6909) );
  BUFX2 U4660 ( .A(n117), .Y(n6910) );
  BUFX2 U4661 ( .A(n151), .Y(n6904) );
  BUFX2 U4662 ( .A(n151), .Y(n6905) );
  BUFX2 U4663 ( .A(n219), .Y(n6894) );
  BUFX2 U4664 ( .A(n219), .Y(n6895) );
  BUFX2 U4665 ( .A(n357), .Y(n6874) );
  BUFX2 U4666 ( .A(n357), .Y(n6875) );
  BUFX2 U4667 ( .A(n391), .Y(n6869) );
  BUFX2 U4668 ( .A(n391), .Y(n6870) );
  BUFX2 U4669 ( .A(n424), .Y(n6864) );
  BUFX2 U4670 ( .A(n424), .Y(n6865) );
  BUFX2 U4671 ( .A(n457), .Y(n6859) );
  BUFX2 U4672 ( .A(n457), .Y(n6860) );
  BUFX2 U4673 ( .A(n490), .Y(n6854) );
  BUFX2 U4674 ( .A(n490), .Y(n6855) );
  BUFX2 U4675 ( .A(n523), .Y(n6849) );
  BUFX2 U4676 ( .A(n523), .Y(n6850) );
  BUFX2 U4677 ( .A(n556), .Y(n6844) );
  BUFX2 U4678 ( .A(n556), .Y(n6845) );
  BUFX2 U4679 ( .A(n589), .Y(n6839) );
  BUFX2 U4680 ( .A(n589), .Y(n6840) );
  BUFX2 U4681 ( .A(n924), .Y(n6789) );
  BUFX2 U4682 ( .A(n924), .Y(n6790) );
  BUFX2 U4683 ( .A(n957), .Y(n6784) );
  BUFX2 U4684 ( .A(n957), .Y(n6785) );
  BUFX2 U4685 ( .A(n990), .Y(n6779) );
  BUFX2 U4686 ( .A(n990), .Y(n6780) );
  BUFX2 U4687 ( .A(n1023), .Y(n6774) );
  BUFX2 U4688 ( .A(n1023), .Y(n6775) );
  BUFX2 U4689 ( .A(n1056), .Y(n6769) );
  BUFX2 U4690 ( .A(n1056), .Y(n6770) );
  BUFX2 U4691 ( .A(n1089), .Y(n6764) );
  BUFX2 U4692 ( .A(n1089), .Y(n6765) );
  BUFX2 U4693 ( .A(n1122), .Y(n6759) );
  BUFX2 U4694 ( .A(n1122), .Y(n6760) );
  BUFX2 U4695 ( .A(n1), .Y(n6927) );
  BUFX2 U4696 ( .A(n1), .Y(n6926) );
  BUFX2 U4697 ( .A(n2096), .Y(n6623) );
  BUFX2 U4698 ( .A(n2164), .Y(n6613) );
  BUFX2 U4699 ( .A(n185), .Y(n6903) );
  BUFX2 U4700 ( .A(n253), .Y(n6893) );
  BUFX2 U4701 ( .A(n624), .Y(n6838) );
  BUFX2 U4702 ( .A(n658), .Y(n6833) );
  BUFX2 U4703 ( .A(n691), .Y(n6828) );
  BUFX2 U4704 ( .A(n724), .Y(n6823) );
  BUFX2 U4705 ( .A(n757), .Y(n6818) );
  BUFX2 U4706 ( .A(n790), .Y(n6813) );
  BUFX2 U4707 ( .A(n823), .Y(n6808) );
  BUFX2 U4708 ( .A(n856), .Y(n6803) );
  BUFX2 U4709 ( .A(n1157), .Y(n6758) );
  BUFX2 U4710 ( .A(n1191), .Y(n6753) );
  BUFX2 U4711 ( .A(n1224), .Y(n6748) );
  BUFX2 U4712 ( .A(n1257), .Y(n6743) );
  BUFX2 U4713 ( .A(n1290), .Y(n6738) );
  BUFX2 U4714 ( .A(n1323), .Y(n6733) );
  BUFX2 U4715 ( .A(n1356), .Y(n6728) );
  BUFX2 U4716 ( .A(n1389), .Y(n6723) );
  BUFX2 U4717 ( .A(n1423), .Y(n6718) );
  BUFX2 U4718 ( .A(n1457), .Y(n6713) );
  BUFX2 U4719 ( .A(n1490), .Y(n6708) );
  BUFX2 U4720 ( .A(n1523), .Y(n6703) );
  BUFX2 U4721 ( .A(n1556), .Y(n6698) );
  BUFX2 U4722 ( .A(n1589), .Y(n6693) );
  BUFX2 U4723 ( .A(n1622), .Y(n6688) );
  BUFX2 U4724 ( .A(n1655), .Y(n6683) );
  BUFX2 U4725 ( .A(n1689), .Y(n6678) );
  BUFX2 U4726 ( .A(n1723), .Y(n6673) );
  BUFX2 U4727 ( .A(n1756), .Y(n6668) );
  BUFX2 U4728 ( .A(n1789), .Y(n6663) );
  BUFX2 U4729 ( .A(n1822), .Y(n6658) );
  BUFX2 U4730 ( .A(n1855), .Y(n6653) );
  BUFX2 U4731 ( .A(n1888), .Y(n6648) );
  BUFX2 U4732 ( .A(n1921), .Y(n6643) );
  BUFX2 U4733 ( .A(n287), .Y(n6888) );
  BUFX2 U4734 ( .A(n321), .Y(n6883) );
  BUFX2 U4735 ( .A(n357), .Y(n6878) );
  BUFX2 U4736 ( .A(n391), .Y(n6873) );
  BUFX2 U4737 ( .A(n424), .Y(n6868) );
  BUFX2 U4738 ( .A(n457), .Y(n6863) );
  BUFX2 U4739 ( .A(n490), .Y(n6858) );
  BUFX2 U4740 ( .A(n523), .Y(n6853) );
  BUFX2 U4741 ( .A(n556), .Y(n6848) );
  BUFX2 U4742 ( .A(n589), .Y(n6843) );
  BUFX2 U4743 ( .A(n2028), .Y(n6633) );
  BUFX2 U4744 ( .A(n2062), .Y(n6628) );
  BUFX2 U4745 ( .A(n2130), .Y(n6618) );
  BUFX2 U4746 ( .A(n82), .Y(n6918) );
  BUFX2 U4747 ( .A(n117), .Y(n6913) );
  BUFX2 U4748 ( .A(n151), .Y(n6908) );
  BUFX2 U4749 ( .A(n219), .Y(n6898) );
  BUFX2 U4750 ( .A(n924), .Y(n6793) );
  BUFX2 U4751 ( .A(n957), .Y(n6788) );
  BUFX2 U4752 ( .A(n990), .Y(n6783) );
  BUFX2 U4753 ( .A(n1023), .Y(n6778) );
  BUFX2 U4754 ( .A(n1056), .Y(n6773) );
  BUFX2 U4755 ( .A(n1089), .Y(n6768) );
  BUFX2 U4756 ( .A(n1122), .Y(n6763) );
  BUFX2 U4757 ( .A(n1), .Y(n6928) );
  BUFX2 U4758 ( .A(n28), .Y(n6923) );
  BUFX2 U4759 ( .A(N13), .Y(n6239) );
  BUFX2 U4760 ( .A(N13), .Y(n6240) );
  BUFX2 U4761 ( .A(N13), .Y(n6241) );
  BUFX2 U4762 ( .A(N13), .Y(n6242) );
  BUFX2 U4763 ( .A(N13), .Y(n6243) );
  BUFX2 U4764 ( .A(N13), .Y(n6244) );
  BUFX2 U4765 ( .A(N13), .Y(n6245) );
  BUFX2 U4766 ( .A(N13), .Y(n6246) );
  BUFX2 U4767 ( .A(N13), .Y(n6247) );
  BUFX2 U4768 ( .A(N14), .Y(n6234) );
  BUFX2 U4769 ( .A(N14), .Y(n6235) );
  BUFX2 U4770 ( .A(N14), .Y(n6236) );
  BUFX2 U4771 ( .A(N14), .Y(n6237) );
  BUFX2 U4772 ( .A(N14), .Y(n6233) );
  BUFX2 U4773 ( .A(N13), .Y(n6238) );
  INVX2 U4774 ( .A(n6231), .Y(n6232) );
  BUFX2 U4775 ( .A(N11), .Y(n6333) );
  BUFX2 U4776 ( .A(N11), .Y(n6332) );
  BUFX2 U4777 ( .A(N11), .Y(n6331) );
  BUFX2 U4778 ( .A(N11), .Y(n6330) );
  BUFX2 U4779 ( .A(N12), .Y(n6269) );
  BUFX2 U4780 ( .A(N12), .Y(n6270) );
  BUFX2 U4781 ( .A(N12), .Y(n6271) );
  BUFX2 U4782 ( .A(N12), .Y(n6272) );
  BUFX2 U4783 ( .A(N12), .Y(n6273) );
  BUFX2 U4784 ( .A(N12), .Y(n6274) );
  BUFX2 U4785 ( .A(N10), .Y(n6448) );
  BUFX2 U4786 ( .A(N10), .Y(n6447) );
  BUFX2 U4787 ( .A(N10), .Y(n6446) );
  BUFX2 U4788 ( .A(N10), .Y(n6445) );
  BUFX2 U4789 ( .A(N10), .Y(n6444) );
  BUFX2 U4790 ( .A(N10), .Y(n6443) );
  BUFX2 U4791 ( .A(N10), .Y(n6442) );
  BUFX2 U4792 ( .A(N10), .Y(n6441) );
  BUFX2 U4793 ( .A(N10), .Y(n6440) );
  BUFX2 U4794 ( .A(N11), .Y(n6329) );
  BUFX2 U4795 ( .A(N12), .Y(n6268) );
  INVX2 U4796 ( .A(RD), .Y(n6939) );
  BUFX2 U4797 ( .A(n7003), .Y(n6604) );
  BUFX2 U4798 ( .A(n6992), .Y(n6549) );
  BUFX2 U4799 ( .A(n6981), .Y(n6494) );
  BUFX2 U4800 ( .A(n6978), .Y(n6479) );
  BUFX2 U4801 ( .A(n6977), .Y(n6474) );
  BUFX2 U4802 ( .A(n6976), .Y(n6469) );
  BUFX2 U4803 ( .A(n6975), .Y(n6464) );
  BUFX2 U4804 ( .A(n6974), .Y(n6459) );
  BUFX2 U4805 ( .A(n6973), .Y(n6454) );
  BUFX2 U4806 ( .A(n6972), .Y(n6449) );
  BUFX2 U4807 ( .A(n7002), .Y(n6599) );
  BUFX2 U4808 ( .A(n7001), .Y(n6594) );
  BUFX2 U4809 ( .A(n7000), .Y(n6589) );
  BUFX2 U4810 ( .A(n6999), .Y(n6584) );
  BUFX2 U4811 ( .A(n6998), .Y(n6579) );
  BUFX2 U4812 ( .A(n6997), .Y(n6574) );
  BUFX2 U4813 ( .A(n6996), .Y(n6569) );
  BUFX2 U4814 ( .A(n6995), .Y(n6564) );
  BUFX2 U4815 ( .A(n6994), .Y(n6559) );
  BUFX2 U4816 ( .A(n6993), .Y(n6554) );
  BUFX2 U4817 ( .A(n6991), .Y(n6544) );
  BUFX2 U4818 ( .A(n6990), .Y(n6539) );
  BUFX2 U4819 ( .A(n6989), .Y(n6534) );
  BUFX2 U4820 ( .A(n6988), .Y(n6529) );
  BUFX2 U4821 ( .A(n6987), .Y(n6524) );
  BUFX2 U4822 ( .A(n6986), .Y(n6519) );
  BUFX2 U4823 ( .A(n6985), .Y(n6514) );
  BUFX2 U4824 ( .A(n6984), .Y(n6509) );
  BUFX2 U4825 ( .A(n6983), .Y(n6504) );
  BUFX2 U4826 ( .A(n6982), .Y(n6499) );
  BUFX2 U4827 ( .A(n6980), .Y(n6489) );
  BUFX2 U4828 ( .A(n6979), .Y(n6484) );
  BUFX2 U4829 ( .A(n7003), .Y(n6605) );
  BUFX2 U4830 ( .A(n6992), .Y(n6550) );
  BUFX2 U4831 ( .A(n6981), .Y(n6495) );
  BUFX2 U4832 ( .A(n6978), .Y(n6480) );
  BUFX2 U4833 ( .A(n6977), .Y(n6475) );
  BUFX2 U4834 ( .A(n6976), .Y(n6470) );
  BUFX2 U4835 ( .A(n6975), .Y(n6465) );
  BUFX2 U4836 ( .A(n6974), .Y(n6460) );
  BUFX2 U4837 ( .A(n6973), .Y(n6455) );
  BUFX2 U4838 ( .A(n6972), .Y(n6450) );
  BUFX2 U4839 ( .A(n7002), .Y(n6600) );
  BUFX2 U4840 ( .A(n7001), .Y(n6595) );
  BUFX2 U4841 ( .A(n7000), .Y(n6590) );
  BUFX2 U4842 ( .A(n6999), .Y(n6585) );
  BUFX2 U4843 ( .A(n6998), .Y(n6580) );
  BUFX2 U4844 ( .A(n6997), .Y(n6575) );
  BUFX2 U4845 ( .A(n6996), .Y(n6570) );
  BUFX2 U4846 ( .A(n6995), .Y(n6565) );
  BUFX2 U4847 ( .A(n6994), .Y(n6560) );
  BUFX2 U4848 ( .A(n6993), .Y(n6555) );
  BUFX2 U4849 ( .A(n6991), .Y(n6545) );
  BUFX2 U4850 ( .A(n6990), .Y(n6540) );
  BUFX2 U4851 ( .A(n6989), .Y(n6535) );
  BUFX2 U4852 ( .A(n6988), .Y(n6530) );
  BUFX2 U4853 ( .A(n6987), .Y(n6525) );
  BUFX2 U4854 ( .A(n6986), .Y(n6520) );
  BUFX2 U4855 ( .A(n6985), .Y(n6515) );
  BUFX2 U4856 ( .A(n6984), .Y(n6510) );
  BUFX2 U4857 ( .A(n6983), .Y(n6505) );
  BUFX2 U4858 ( .A(n6982), .Y(n6500) );
  BUFX2 U4859 ( .A(n6980), .Y(n6490) );
  BUFX2 U4860 ( .A(n6979), .Y(n6485) );
  BUFX2 U4861 ( .A(n7003), .Y(n6606) );
  BUFX2 U4862 ( .A(n6992), .Y(n6551) );
  BUFX2 U4863 ( .A(n6981), .Y(n6496) );
  BUFX2 U4864 ( .A(n6978), .Y(n6481) );
  BUFX2 U4865 ( .A(n6977), .Y(n6476) );
  BUFX2 U4866 ( .A(n6976), .Y(n6471) );
  BUFX2 U4867 ( .A(n6975), .Y(n6466) );
  BUFX2 U4868 ( .A(n6974), .Y(n6461) );
  BUFX2 U4869 ( .A(n6973), .Y(n6456) );
  BUFX2 U4870 ( .A(n6972), .Y(n6451) );
  BUFX2 U4871 ( .A(n7002), .Y(n6601) );
  BUFX2 U4872 ( .A(n7001), .Y(n6596) );
  BUFX2 U4873 ( .A(n7000), .Y(n6591) );
  BUFX2 U4874 ( .A(n6999), .Y(n6586) );
  BUFX2 U4875 ( .A(n6998), .Y(n6581) );
  BUFX2 U4876 ( .A(n6997), .Y(n6576) );
  BUFX2 U4877 ( .A(n6996), .Y(n6571) );
  BUFX2 U4878 ( .A(n6995), .Y(n6566) );
  BUFX2 U4879 ( .A(n6994), .Y(n6561) );
  BUFX2 U4880 ( .A(n6993), .Y(n6556) );
  BUFX2 U4881 ( .A(n6991), .Y(n6546) );
  BUFX2 U4882 ( .A(n6990), .Y(n6541) );
  BUFX2 U4883 ( .A(n6989), .Y(n6536) );
  BUFX2 U4884 ( .A(n6988), .Y(n6531) );
  BUFX2 U4885 ( .A(n6987), .Y(n6526) );
  BUFX2 U4886 ( .A(n6986), .Y(n6521) );
  BUFX2 U4887 ( .A(n6985), .Y(n6516) );
  BUFX2 U4888 ( .A(n6984), .Y(n6511) );
  BUFX2 U4889 ( .A(n6983), .Y(n6506) );
  BUFX2 U4890 ( .A(n6982), .Y(n6501) );
  BUFX2 U4891 ( .A(n6980), .Y(n6491) );
  BUFX2 U4892 ( .A(n6979), .Y(n6486) );
  BUFX2 U4893 ( .A(n7003), .Y(n6607) );
  BUFX2 U4894 ( .A(n6992), .Y(n6552) );
  BUFX2 U4895 ( .A(n6981), .Y(n6497) );
  BUFX2 U4896 ( .A(n6978), .Y(n6482) );
  BUFX2 U4897 ( .A(n6977), .Y(n6477) );
  BUFX2 U4898 ( .A(n6976), .Y(n6472) );
  BUFX2 U4899 ( .A(n6975), .Y(n6467) );
  BUFX2 U4900 ( .A(n6974), .Y(n6462) );
  BUFX2 U4901 ( .A(n6973), .Y(n6457) );
  BUFX2 U4902 ( .A(n6972), .Y(n6452) );
  BUFX2 U4903 ( .A(n7002), .Y(n6602) );
  BUFX2 U4904 ( .A(n7001), .Y(n6597) );
  BUFX2 U4905 ( .A(n7000), .Y(n6592) );
  BUFX2 U4906 ( .A(n6999), .Y(n6587) );
  BUFX2 U4907 ( .A(n6998), .Y(n6582) );
  BUFX2 U4908 ( .A(n6997), .Y(n6577) );
  BUFX2 U4909 ( .A(n6996), .Y(n6572) );
  BUFX2 U4910 ( .A(n6995), .Y(n6567) );
  BUFX2 U4911 ( .A(n6994), .Y(n6562) );
  BUFX2 U4912 ( .A(n6993), .Y(n6557) );
  BUFX2 U4913 ( .A(n6991), .Y(n6547) );
  BUFX2 U4914 ( .A(n6990), .Y(n6542) );
  BUFX2 U4915 ( .A(n6989), .Y(n6537) );
  BUFX2 U4916 ( .A(n6988), .Y(n6532) );
  BUFX2 U4917 ( .A(n6987), .Y(n6527) );
  BUFX2 U4918 ( .A(n6986), .Y(n6522) );
  BUFX2 U4919 ( .A(n6985), .Y(n6517) );
  BUFX2 U4920 ( .A(n6984), .Y(n6512) );
  BUFX2 U4921 ( .A(n6983), .Y(n6507) );
  BUFX2 U4922 ( .A(n6982), .Y(n6502) );
  BUFX2 U4923 ( .A(n6980), .Y(n6492) );
  BUFX2 U4924 ( .A(n6979), .Y(n6487) );
  BUFX2 U4925 ( .A(n7003), .Y(n6608) );
  BUFX2 U4926 ( .A(n6992), .Y(n6553) );
  BUFX2 U4927 ( .A(n6972), .Y(n6453) );
  BUFX2 U4928 ( .A(n7002), .Y(n6603) );
  BUFX2 U4929 ( .A(n7001), .Y(n6598) );
  BUFX2 U4930 ( .A(n7000), .Y(n6593) );
  BUFX2 U4931 ( .A(n6999), .Y(n6588) );
  BUFX2 U4932 ( .A(n6998), .Y(n6583) );
  BUFX2 U4933 ( .A(n6997), .Y(n6578) );
  BUFX2 U4934 ( .A(n6995), .Y(n6568) );
  BUFX2 U4935 ( .A(n6994), .Y(n6563) );
  BUFX2 U4936 ( .A(n6993), .Y(n6558) );
  BUFX2 U4937 ( .A(n6991), .Y(n6548) );
  BUFX2 U4938 ( .A(n6990), .Y(n6543) );
  BUFX2 U4939 ( .A(n6981), .Y(n6498) );
  BUFX2 U4940 ( .A(n6978), .Y(n6483) );
  BUFX2 U4941 ( .A(n6977), .Y(n6478) );
  BUFX2 U4942 ( .A(n6976), .Y(n6473) );
  BUFX2 U4943 ( .A(n6975), .Y(n6468) );
  BUFX2 U4944 ( .A(n6974), .Y(n6463) );
  BUFX2 U4945 ( .A(n6973), .Y(n6458) );
  BUFX2 U4946 ( .A(n6996), .Y(n6573) );
  BUFX2 U4947 ( .A(n6989), .Y(n6538) );
  BUFX2 U4948 ( .A(n6988), .Y(n6533) );
  BUFX2 U4949 ( .A(n6987), .Y(n6528) );
  BUFX2 U4950 ( .A(n6986), .Y(n6523) );
  BUFX2 U4951 ( .A(n6985), .Y(n6518) );
  BUFX2 U4952 ( .A(n6984), .Y(n6513) );
  BUFX2 U4953 ( .A(n6983), .Y(n6508) );
  BUFX2 U4954 ( .A(n6982), .Y(n6503) );
  BUFX2 U4955 ( .A(n6980), .Y(n6493) );
  BUFX2 U4956 ( .A(n6979), .Y(n6488) );
  INVX2 U4957 ( .A(N15), .Y(n6231) );
  MUX2X1 U4958 ( .B(n116), .A(n150), .S(n6289), .Y(n115) );
  MUX2X1 U4959 ( .B(n218), .A(n252), .S(n6289), .Y(n184) );
  MUX2X1 U4960 ( .B(n320), .A(n356), .S(n6289), .Y(n286) );
  MUX2X1 U4961 ( .B(n623), .A(n657), .S(n6289), .Y(n390) );
  MUX2X1 U4962 ( .B(n1190), .A(n1456), .S(n6238), .Y(n923) );
  MUX2X1 U4963 ( .B(n1956), .A(n1959), .S(n6289), .Y(n1722) );
  MUX2X1 U4964 ( .B(n2026), .A(n2027), .S(n6290), .Y(n2025) );
  MUX2X1 U4965 ( .B(n2221), .A(n2222), .S(n6290), .Y(n2218) );
  MUX2X1 U4966 ( .B(n2224), .A(n2225), .S(n6290), .Y(n2223) );
  MUX2X1 U4967 ( .B(n2227), .A(n2228), .S(n6238), .Y(n2226) );
  MUX2X1 U4968 ( .B(n2230), .A(n2231), .S(n6290), .Y(n2229) );
  MUX2X1 U4969 ( .B(n2233), .A(n2234), .S(n6290), .Y(n2232) );
  MUX2X1 U4970 ( .B(n2236), .A(n2237), .S(n6290), .Y(n2235) );
  MUX2X1 U4971 ( .B(n2239), .A(n2240), .S(n6290), .Y(n2238) );
  MUX2X1 U4972 ( .B(n2242), .A(n2243), .S(n6238), .Y(n2241) );
  MUX2X1 U4973 ( .B(n2245), .A(n2246), .S(n6290), .Y(n2244) );
  MUX2X1 U4974 ( .B(n2248), .A(n2249), .S(n6290), .Y(n2247) );
  MUX2X1 U4975 ( .B(n2251), .A(n2252), .S(n6290), .Y(n2250) );
  MUX2X1 U4976 ( .B(n2254), .A(n2255), .S(n6290), .Y(n2253) );
  MUX2X1 U4977 ( .B(n2257), .A(n2258), .S(n6238), .Y(n2256) );
  MUX2X1 U4978 ( .B(n2259), .A(n2260), .S(N15), .Y(N112) );
  MUX2X1 U4979 ( .B(n2262), .A(n2263), .S(n6290), .Y(n2261) );
  MUX2X1 U4980 ( .B(n2265), .A(n2266), .S(n6290), .Y(n2264) );
  MUX2X1 U4981 ( .B(n2268), .A(n2269), .S(n6291), .Y(n2267) );
  MUX2X1 U4982 ( .B(n2271), .A(n2272), .S(n6291), .Y(n2270) );
  MUX2X1 U4983 ( .B(n2274), .A(n2275), .S(n6238), .Y(n2273) );
  MUX2X1 U4984 ( .B(n2277), .A(n2278), .S(n6291), .Y(n2276) );
  MUX2X1 U4985 ( .B(n2280), .A(n2281), .S(n6291), .Y(n2279) );
  MUX2X1 U4986 ( .B(n2283), .A(n2284), .S(n6291), .Y(n2282) );
  MUX2X1 U4987 ( .B(n4334), .A(n4335), .S(n6291), .Y(n2285) );
  MUX2X1 U4988 ( .B(n4337), .A(n4338), .S(n6238), .Y(n4336) );
  MUX2X1 U4989 ( .B(n4340), .A(n4341), .S(n6291), .Y(n4339) );
  MUX2X1 U4990 ( .B(n4343), .A(n4344), .S(n6291), .Y(n4342) );
  MUX2X1 U4991 ( .B(n4346), .A(n4347), .S(n6291), .Y(n4345) );
  MUX2X1 U4992 ( .B(n4349), .A(n4350), .S(n6291), .Y(n4348) );
  MUX2X1 U4993 ( .B(n4352), .A(n4353), .S(n6238), .Y(n4351) );
  MUX2X1 U4994 ( .B(n4355), .A(n4356), .S(n6291), .Y(n4354) );
  MUX2X1 U4995 ( .B(n4358), .A(n4359), .S(n6291), .Y(n4357) );
  MUX2X1 U4996 ( .B(n4361), .A(n4362), .S(n6291), .Y(n4360) );
  MUX2X1 U4997 ( .B(n4364), .A(n4365), .S(n6292), .Y(n4363) );
  MUX2X1 U4998 ( .B(n4367), .A(n4368), .S(n6238), .Y(n4366) );
  MUX2X1 U4999 ( .B(n4369), .A(n4370), .S(N15), .Y(N111) );
  MUX2X1 U5000 ( .B(n4372), .A(n4373), .S(n6292), .Y(n4371) );
  MUX2X1 U5001 ( .B(n4375), .A(n4376), .S(n6292), .Y(n4374) );
  MUX2X1 U5002 ( .B(n4378), .A(n4379), .S(n6292), .Y(n4377) );
  MUX2X1 U5003 ( .B(n4381), .A(n4382), .S(n6292), .Y(n4380) );
  MUX2X1 U5004 ( .B(n4384), .A(n4385), .S(n6238), .Y(n4383) );
  MUX2X1 U5005 ( .B(n4387), .A(n4388), .S(n6292), .Y(n4386) );
  MUX2X1 U5006 ( .B(n4390), .A(n4391), .S(n6292), .Y(n4389) );
  MUX2X1 U5007 ( .B(n4393), .A(n4394), .S(n6292), .Y(n4392) );
  MUX2X1 U5008 ( .B(n4396), .A(n4397), .S(n6292), .Y(n4395) );
  MUX2X1 U5009 ( .B(n4399), .A(n4400), .S(n6238), .Y(n4398) );
  MUX2X1 U5010 ( .B(n4402), .A(n4403), .S(n6292), .Y(n4401) );
  MUX2X1 U5011 ( .B(n4405), .A(n4406), .S(n6292), .Y(n4404) );
  MUX2X1 U5012 ( .B(n4408), .A(n4409), .S(n6292), .Y(n4407) );
  MUX2X1 U5013 ( .B(n4411), .A(n4412), .S(n6292), .Y(n4410) );
  MUX2X1 U5014 ( .B(n4414), .A(n4415), .S(n6238), .Y(n4413) );
  MUX2X1 U5015 ( .B(n4417), .A(n4418), .S(n6293), .Y(n4416) );
  MUX2X1 U5016 ( .B(n4420), .A(n4421), .S(n6293), .Y(n4419) );
  MUX2X1 U5017 ( .B(n4423), .A(n4424), .S(n6293), .Y(n4422) );
  MUX2X1 U5018 ( .B(n4426), .A(n4427), .S(n6293), .Y(n4425) );
  MUX2X1 U5019 ( .B(n4429), .A(n4430), .S(n6239), .Y(n4428) );
  MUX2X1 U5020 ( .B(n4431), .A(n4432), .S(N15), .Y(N110) );
  MUX2X1 U5021 ( .B(n4434), .A(n4435), .S(n6293), .Y(n4433) );
  MUX2X1 U5022 ( .B(n4437), .A(n4438), .S(n6293), .Y(n4436) );
  MUX2X1 U5023 ( .B(n4440), .A(n4441), .S(n6293), .Y(n4439) );
  MUX2X1 U5024 ( .B(n4443), .A(n4444), .S(n6293), .Y(n4442) );
  MUX2X1 U5025 ( .B(n4446), .A(n4447), .S(n6239), .Y(n4445) );
  MUX2X1 U5026 ( .B(n4449), .A(n4450), .S(n6293), .Y(n4448) );
  MUX2X1 U5027 ( .B(n4452), .A(n4453), .S(n6293), .Y(n4451) );
  MUX2X1 U5028 ( .B(n4455), .A(n4456), .S(n6293), .Y(n4454) );
  MUX2X1 U5029 ( .B(n4458), .A(n4459), .S(n6293), .Y(n4457) );
  MUX2X1 U5030 ( .B(n4461), .A(n4462), .S(n6239), .Y(n4460) );
  MUX2X1 U5031 ( .B(n4464), .A(n4465), .S(n6293), .Y(n4463) );
  MUX2X1 U5032 ( .B(n4467), .A(n4468), .S(n6294), .Y(n4466) );
  MUX2X1 U5033 ( .B(n4470), .A(n4471), .S(n6294), .Y(n4469) );
  MUX2X1 U5034 ( .B(n4473), .A(n4474), .S(n6294), .Y(n4472) );
  MUX2X1 U5035 ( .B(n4476), .A(n4477), .S(n6239), .Y(n4475) );
  MUX2X1 U5036 ( .B(n4479), .A(n4480), .S(n6294), .Y(n4478) );
  MUX2X1 U5037 ( .B(n4482), .A(n4483), .S(n6294), .Y(n4481) );
  MUX2X1 U5038 ( .B(n4485), .A(n4486), .S(n6294), .Y(n4484) );
  MUX2X1 U5039 ( .B(n4488), .A(n4489), .S(n6294), .Y(n4487) );
  MUX2X1 U5040 ( .B(n4491), .A(n4492), .S(n6239), .Y(n4490) );
  MUX2X1 U5041 ( .B(n4493), .A(n4494), .S(N15), .Y(N109) );
  MUX2X1 U5042 ( .B(n4496), .A(n4497), .S(n6294), .Y(n4495) );
  MUX2X1 U5043 ( .B(n4499), .A(n4500), .S(n6294), .Y(n4498) );
  MUX2X1 U5044 ( .B(n4502), .A(n4503), .S(n6294), .Y(n4501) );
  MUX2X1 U5045 ( .B(n4505), .A(n4506), .S(n6294), .Y(n4504) );
  MUX2X1 U5046 ( .B(n4508), .A(n4509), .S(n6239), .Y(n4507) );
  MUX2X1 U5047 ( .B(n4511), .A(n4512), .S(n6294), .Y(n4510) );
  MUX2X1 U5048 ( .B(n4514), .A(n4515), .S(n6294), .Y(n4513) );
  MUX2X1 U5049 ( .B(n4517), .A(n4518), .S(n6295), .Y(n4516) );
  MUX2X1 U5050 ( .B(n4520), .A(n4521), .S(n6295), .Y(n4519) );
  MUX2X1 U5051 ( .B(n4523), .A(n4524), .S(n6239), .Y(n4522) );
  MUX2X1 U5052 ( .B(n4526), .A(n4527), .S(n6295), .Y(n4525) );
  MUX2X1 U5053 ( .B(n4529), .A(n4530), .S(n6295), .Y(n4528) );
  MUX2X1 U5054 ( .B(n4532), .A(n4533), .S(n6295), .Y(n4531) );
  MUX2X1 U5055 ( .B(n4535), .A(n4536), .S(n6295), .Y(n4534) );
  MUX2X1 U5056 ( .B(n4538), .A(n4539), .S(n6239), .Y(n4537) );
  MUX2X1 U5057 ( .B(n4541), .A(n4542), .S(n6295), .Y(n4540) );
  MUX2X1 U5058 ( .B(n4544), .A(n4545), .S(n6295), .Y(n4543) );
  MUX2X1 U5059 ( .B(n4547), .A(n4548), .S(n6295), .Y(n4546) );
  MUX2X1 U5060 ( .B(n4550), .A(n4551), .S(n6295), .Y(n4549) );
  MUX2X1 U5061 ( .B(n4553), .A(n4554), .S(n6239), .Y(n4552) );
  MUX2X1 U5062 ( .B(n4555), .A(n4556), .S(N15), .Y(N108) );
  MUX2X1 U5063 ( .B(n4558), .A(n4559), .S(n6295), .Y(n4557) );
  MUX2X1 U5064 ( .B(n4561), .A(n4562), .S(n6295), .Y(n4560) );
  MUX2X1 U5065 ( .B(n4564), .A(n4565), .S(n6295), .Y(n4563) );
  MUX2X1 U5066 ( .B(n4567), .A(n4568), .S(n6296), .Y(n4566) );
  MUX2X1 U5067 ( .B(n4570), .A(n4571), .S(n6239), .Y(n4569) );
  MUX2X1 U5068 ( .B(n4573), .A(n4574), .S(n6296), .Y(n4572) );
  MUX2X1 U5069 ( .B(n4576), .A(n4577), .S(n6296), .Y(n4575) );
  MUX2X1 U5070 ( .B(n4579), .A(n4580), .S(n6296), .Y(n4578) );
  MUX2X1 U5071 ( .B(n4582), .A(n4583), .S(n6296), .Y(n4581) );
  MUX2X1 U5072 ( .B(n4585), .A(n4586), .S(n6239), .Y(n4584) );
  MUX2X1 U5073 ( .B(n4588), .A(n4589), .S(n6296), .Y(n4587) );
  MUX2X1 U5074 ( .B(n4591), .A(n4592), .S(n6296), .Y(n4590) );
  MUX2X1 U5075 ( .B(n4594), .A(n4595), .S(n6296), .Y(n4593) );
  MUX2X1 U5076 ( .B(n4597), .A(n4598), .S(n6296), .Y(n4596) );
  MUX2X1 U5077 ( .B(n4600), .A(n4601), .S(n6239), .Y(n4599) );
  MUX2X1 U5078 ( .B(n4603), .A(n4604), .S(n6296), .Y(n4602) );
  MUX2X1 U5079 ( .B(n4606), .A(n4607), .S(n6296), .Y(n4605) );
  MUX2X1 U5080 ( .B(n4609), .A(n4610), .S(n6296), .Y(n4608) );
  MUX2X1 U5081 ( .B(n4612), .A(n4613), .S(n6296), .Y(n4611) );
  MUX2X1 U5082 ( .B(n4615), .A(n4616), .S(n6239), .Y(n4614) );
  MUX2X1 U5083 ( .B(n4617), .A(n4618), .S(N15), .Y(N107) );
  MUX2X1 U5084 ( .B(n4620), .A(n4621), .S(n6297), .Y(n4619) );
  MUX2X1 U5085 ( .B(n4623), .A(n4624), .S(n6297), .Y(n4622) );
  MUX2X1 U5086 ( .B(n4626), .A(n4627), .S(n6297), .Y(n4625) );
  MUX2X1 U5087 ( .B(n4629), .A(n4630), .S(n6297), .Y(n4628) );
  MUX2X1 U5088 ( .B(n4632), .A(n4633), .S(n6240), .Y(n4631) );
  MUX2X1 U5089 ( .B(n4635), .A(n4636), .S(n6297), .Y(n4634) );
  MUX2X1 U5090 ( .B(n4638), .A(n4639), .S(n6297), .Y(n4637) );
  MUX2X1 U5091 ( .B(n4641), .A(n4642), .S(n6297), .Y(n4640) );
  MUX2X1 U5092 ( .B(n4644), .A(n4645), .S(n6297), .Y(n4643) );
  MUX2X1 U5093 ( .B(n4647), .A(n4648), .S(n6240), .Y(n4646) );
  MUX2X1 U5094 ( .B(n4650), .A(n4651), .S(n6297), .Y(n4649) );
  MUX2X1 U5095 ( .B(n4653), .A(n4654), .S(n6297), .Y(n4652) );
  MUX2X1 U5096 ( .B(n4656), .A(n4657), .S(n6297), .Y(n4655) );
  MUX2X1 U5097 ( .B(n4659), .A(n4660), .S(n6297), .Y(n4658) );
  MUX2X1 U5098 ( .B(n4662), .A(n4663), .S(n6240), .Y(n4661) );
  MUX2X1 U5099 ( .B(n4665), .A(n4666), .S(n6297), .Y(n4664) );
  MUX2X1 U5100 ( .B(n4668), .A(n4669), .S(n6298), .Y(n4667) );
  MUX2X1 U5101 ( .B(n4671), .A(n4672), .S(n6298), .Y(n4670) );
  MUX2X1 U5102 ( .B(n4674), .A(n4675), .S(n6298), .Y(n4673) );
  MUX2X1 U5103 ( .B(n4677), .A(n4678), .S(n6240), .Y(n4676) );
  MUX2X1 U5104 ( .B(n4679), .A(n4680), .S(n6232), .Y(N106) );
  MUX2X1 U5105 ( .B(n4682), .A(n4683), .S(n6298), .Y(n4681) );
  MUX2X1 U5106 ( .B(n4685), .A(n4686), .S(n6298), .Y(n4684) );
  MUX2X1 U5107 ( .B(n4688), .A(n4689), .S(n6298), .Y(n4687) );
  MUX2X1 U5108 ( .B(n4691), .A(n4692), .S(n6298), .Y(n4690) );
  MUX2X1 U5109 ( .B(n4694), .A(n4695), .S(n6240), .Y(n4693) );
  MUX2X1 U5110 ( .B(n4697), .A(n4698), .S(n6298), .Y(n4696) );
  MUX2X1 U5111 ( .B(n4700), .A(n4701), .S(n6298), .Y(n4699) );
  MUX2X1 U5112 ( .B(n4703), .A(n4704), .S(n6298), .Y(n4702) );
  MUX2X1 U5113 ( .B(n4706), .A(n4707), .S(n6298), .Y(n4705) );
  MUX2X1 U5114 ( .B(n4709), .A(n4710), .S(n6240), .Y(n4708) );
  MUX2X1 U5115 ( .B(n4712), .A(n4713), .S(n6298), .Y(n4711) );
  MUX2X1 U5116 ( .B(n4715), .A(n4716), .S(n6298), .Y(n4714) );
  MUX2X1 U5117 ( .B(n4718), .A(n4719), .S(n6299), .Y(n4717) );
  MUX2X1 U5118 ( .B(n4721), .A(n4722), .S(n6299), .Y(n4720) );
  MUX2X1 U5119 ( .B(n4724), .A(n4725), .S(n6240), .Y(n4723) );
  MUX2X1 U5120 ( .B(n4727), .A(n4728), .S(n6299), .Y(n4726) );
  MUX2X1 U5121 ( .B(n4730), .A(n4731), .S(n6299), .Y(n4729) );
  MUX2X1 U5122 ( .B(n4733), .A(n4734), .S(n6299), .Y(n4732) );
  MUX2X1 U5123 ( .B(n4736), .A(n4737), .S(n6299), .Y(n4735) );
  MUX2X1 U5124 ( .B(n4739), .A(n4740), .S(n6240), .Y(n4738) );
  MUX2X1 U5125 ( .B(n4741), .A(n4742), .S(n6232), .Y(N105) );
  MUX2X1 U5126 ( .B(n4744), .A(n4745), .S(n6299), .Y(n4743) );
  MUX2X1 U5127 ( .B(n4747), .A(n4748), .S(n6299), .Y(n4746) );
  MUX2X1 U5128 ( .B(n4750), .A(n4751), .S(n6299), .Y(n4749) );
  MUX2X1 U5129 ( .B(n4753), .A(n4754), .S(n6299), .Y(n4752) );
  MUX2X1 U5130 ( .B(n4756), .A(n4757), .S(n6240), .Y(n4755) );
  MUX2X1 U5131 ( .B(n4759), .A(n4760), .S(n6299), .Y(n4758) );
  MUX2X1 U5132 ( .B(n4762), .A(n4763), .S(n6299), .Y(n4761) );
  MUX2X1 U5133 ( .B(n4765), .A(n4766), .S(n6299), .Y(n4764) );
  MUX2X1 U5134 ( .B(n4768), .A(n4769), .S(n6300), .Y(n4767) );
  MUX2X1 U5135 ( .B(n4771), .A(n4772), .S(n6240), .Y(n4770) );
  MUX2X1 U5136 ( .B(n4774), .A(n4775), .S(n6300), .Y(n4773) );
  MUX2X1 U5137 ( .B(n4777), .A(n4778), .S(n6300), .Y(n4776) );
  MUX2X1 U5138 ( .B(n4780), .A(n4781), .S(n6300), .Y(n4779) );
  MUX2X1 U5139 ( .B(n4783), .A(n4784), .S(n6300), .Y(n4782) );
  MUX2X1 U5140 ( .B(n4786), .A(n4787), .S(n6240), .Y(n4785) );
  MUX2X1 U5141 ( .B(n4789), .A(n4790), .S(n6300), .Y(n4788) );
  MUX2X1 U5142 ( .B(n4792), .A(n4793), .S(n6300), .Y(n4791) );
  MUX2X1 U5143 ( .B(n4795), .A(n4796), .S(n6300), .Y(n4794) );
  MUX2X1 U5144 ( .B(n4798), .A(n4799), .S(n6300), .Y(n4797) );
  MUX2X1 U5145 ( .B(n4801), .A(n4802), .S(n6240), .Y(n4800) );
  MUX2X1 U5146 ( .B(n4803), .A(n4804), .S(n6232), .Y(N104) );
  MUX2X1 U5147 ( .B(n4806), .A(n4807), .S(n6300), .Y(n4805) );
  MUX2X1 U5148 ( .B(n4809), .A(n4810), .S(n6300), .Y(n4808) );
  MUX2X1 U5149 ( .B(n4812), .A(n4813), .S(n6300), .Y(n4811) );
  MUX2X1 U5150 ( .B(n4815), .A(n4816), .S(n6300), .Y(n4814) );
  MUX2X1 U5151 ( .B(n4818), .A(n4819), .S(n6240), .Y(n4817) );
  MUX2X1 U5152 ( .B(n4821), .A(n4822), .S(n6301), .Y(n4820) );
  MUX2X1 U5153 ( .B(n4824), .A(n4825), .S(n6301), .Y(n4823) );
  MUX2X1 U5154 ( .B(n4827), .A(n4828), .S(n6301), .Y(n4826) );
  MUX2X1 U5155 ( .B(n4830), .A(n4831), .S(n6301), .Y(n4829) );
  MUX2X1 U5156 ( .B(n4833), .A(n4834), .S(n6241), .Y(n4832) );
  MUX2X1 U5157 ( .B(n4836), .A(n4837), .S(n6301), .Y(n4835) );
  MUX2X1 U5158 ( .B(n4839), .A(n4840), .S(n6301), .Y(n4838) );
  MUX2X1 U5159 ( .B(n4842), .A(n4843), .S(n6301), .Y(n4841) );
  MUX2X1 U5160 ( .B(n4845), .A(n4846), .S(n6301), .Y(n4844) );
  MUX2X1 U5161 ( .B(n4848), .A(n4849), .S(n6241), .Y(n4847) );
  MUX2X1 U5162 ( .B(n4851), .A(n4852), .S(n6301), .Y(n4850) );
  MUX2X1 U5163 ( .B(n4854), .A(n4855), .S(n6301), .Y(n4853) );
  MUX2X1 U5164 ( .B(n4857), .A(n4858), .S(n6301), .Y(n4856) );
  MUX2X1 U5165 ( .B(n4860), .A(n4861), .S(n6301), .Y(n4859) );
  MUX2X1 U5166 ( .B(n4863), .A(n4864), .S(n6241), .Y(n4862) );
  MUX2X1 U5167 ( .B(n4865), .A(n4866), .S(n6232), .Y(N103) );
  MUX2X1 U5168 ( .B(n4868), .A(n4869), .S(n6301), .Y(n4867) );
  MUX2X1 U5169 ( .B(n4871), .A(n4872), .S(n6302), .Y(n4870) );
  MUX2X1 U5170 ( .B(n4874), .A(n4875), .S(n6302), .Y(n4873) );
  MUX2X1 U5171 ( .B(n4877), .A(n4878), .S(n6302), .Y(n4876) );
  MUX2X1 U5172 ( .B(n4880), .A(n4881), .S(n6241), .Y(n4879) );
  MUX2X1 U5173 ( .B(n4883), .A(n4884), .S(n6302), .Y(n4882) );
  MUX2X1 U5174 ( .B(n4886), .A(n4887), .S(n6302), .Y(n4885) );
  MUX2X1 U5175 ( .B(n4889), .A(n4890), .S(n6302), .Y(n4888) );
  MUX2X1 U5176 ( .B(n4892), .A(n4893), .S(n6302), .Y(n4891) );
  MUX2X1 U5177 ( .B(n4895), .A(n4896), .S(n6241), .Y(n4894) );
  MUX2X1 U5178 ( .B(n4898), .A(n4899), .S(n6302), .Y(n4897) );
  MUX2X1 U5179 ( .B(n4901), .A(n4902), .S(n6302), .Y(n4900) );
  MUX2X1 U5180 ( .B(n4904), .A(n4905), .S(n6302), .Y(n4903) );
  MUX2X1 U5181 ( .B(n4907), .A(n4908), .S(n6302), .Y(n4906) );
  MUX2X1 U5182 ( .B(n4910), .A(n4911), .S(n6241), .Y(n4909) );
  MUX2X1 U5183 ( .B(n4913), .A(n4914), .S(n6302), .Y(n4912) );
  MUX2X1 U5184 ( .B(n4916), .A(n4917), .S(n6302), .Y(n4915) );
  MUX2X1 U5185 ( .B(n4919), .A(n4920), .S(n6303), .Y(n4918) );
  MUX2X1 U5186 ( .B(n4922), .A(n4923), .S(n6303), .Y(n4921) );
  MUX2X1 U5187 ( .B(n4925), .A(n4926), .S(n6241), .Y(n4924) );
  MUX2X1 U5188 ( .B(n4927), .A(n4928), .S(n6232), .Y(N102) );
  MUX2X1 U5189 ( .B(n4930), .A(n4931), .S(n6303), .Y(n4929) );
  MUX2X1 U5190 ( .B(n4933), .A(n4934), .S(n6303), .Y(n4932) );
  MUX2X1 U5191 ( .B(n4936), .A(n4937), .S(n6303), .Y(n4935) );
  MUX2X1 U5192 ( .B(n4939), .A(n4940), .S(n6303), .Y(n4938) );
  MUX2X1 U5193 ( .B(n4942), .A(n4943), .S(n6241), .Y(n4941) );
  MUX2X1 U5194 ( .B(n4945), .A(n4946), .S(n6303), .Y(n4944) );
  MUX2X1 U5195 ( .B(n4948), .A(n4949), .S(n6303), .Y(n4947) );
  MUX2X1 U5196 ( .B(n4951), .A(n4952), .S(n6303), .Y(n4950) );
  MUX2X1 U5197 ( .B(n4954), .A(n4955), .S(n6303), .Y(n4953) );
  MUX2X1 U5198 ( .B(n4957), .A(n4958), .S(n6241), .Y(n4956) );
  MUX2X1 U5199 ( .B(n4960), .A(n4961), .S(n6303), .Y(n4959) );
  MUX2X1 U5200 ( .B(n4963), .A(n4964), .S(n6303), .Y(n4962) );
  MUX2X1 U5201 ( .B(n4966), .A(n4967), .S(n6303), .Y(n4965) );
  MUX2X1 U5202 ( .B(n4969), .A(n4970), .S(n6304), .Y(n4968) );
  MUX2X1 U5203 ( .B(n4972), .A(n4973), .S(n6241), .Y(n4971) );
  MUX2X1 U5204 ( .B(n4975), .A(n4976), .S(n6304), .Y(n4974) );
  MUX2X1 U5205 ( .B(n4978), .A(n4979), .S(n6304), .Y(n4977) );
  MUX2X1 U5206 ( .B(n4981), .A(n4982), .S(n6304), .Y(n4980) );
  MUX2X1 U5207 ( .B(n4984), .A(n4985), .S(n6304), .Y(n4983) );
  MUX2X1 U5208 ( .B(n4987), .A(n4988), .S(n6241), .Y(n4986) );
  MUX2X1 U5209 ( .B(n4989), .A(n4990), .S(n6232), .Y(N101) );
  MUX2X1 U5210 ( .B(n4992), .A(n4993), .S(n6304), .Y(n4991) );
  MUX2X1 U5211 ( .B(n4995), .A(n4996), .S(n6304), .Y(n4994) );
  MUX2X1 U5212 ( .B(n4998), .A(n4999), .S(n6304), .Y(n4997) );
  MUX2X1 U5213 ( .B(n5001), .A(n5002), .S(n6304), .Y(n5000) );
  MUX2X1 U5214 ( .B(n5004), .A(n5005), .S(n6241), .Y(n5003) );
  MUX2X1 U5215 ( .B(n5007), .A(n5008), .S(n6304), .Y(n5006) );
  MUX2X1 U5216 ( .B(n5010), .A(n5011), .S(n6304), .Y(n5009) );
  MUX2X1 U5217 ( .B(n5013), .A(n5014), .S(n6304), .Y(n5012) );
  MUX2X1 U5218 ( .B(n5016), .A(n5017), .S(n6304), .Y(n5015) );
  MUX2X1 U5219 ( .B(n5019), .A(n5020), .S(n6241), .Y(n5018) );
  MUX2X1 U5220 ( .B(n5022), .A(n5023), .S(n6305), .Y(n5021) );
  MUX2X1 U5221 ( .B(n5025), .A(n5026), .S(n6305), .Y(n5024) );
  MUX2X1 U5222 ( .B(n5028), .A(n5029), .S(n6305), .Y(n5027) );
  MUX2X1 U5223 ( .B(n5031), .A(n5032), .S(n6305), .Y(n5030) );
  MUX2X1 U5224 ( .B(n5034), .A(n5035), .S(n6242), .Y(n5033) );
  MUX2X1 U5225 ( .B(n5037), .A(n5038), .S(n6305), .Y(n5036) );
  MUX2X1 U5226 ( .B(n5040), .A(n5041), .S(n6305), .Y(n5039) );
  MUX2X1 U5227 ( .B(n5043), .A(n5044), .S(n6305), .Y(n5042) );
  MUX2X1 U5228 ( .B(n5046), .A(n5047), .S(n6305), .Y(n5045) );
  MUX2X1 U5229 ( .B(n5049), .A(n5050), .S(n6242), .Y(n5048) );
  MUX2X1 U5230 ( .B(n5051), .A(n5052), .S(n6232), .Y(N100) );
  MUX2X1 U5231 ( .B(n5054), .A(n5055), .S(n6305), .Y(n5053) );
  MUX2X1 U5232 ( .B(n5057), .A(n5058), .S(n6305), .Y(n5056) );
  MUX2X1 U5233 ( .B(n5060), .A(n5061), .S(n6305), .Y(n5059) );
  MUX2X1 U5234 ( .B(n5063), .A(n5064), .S(n6305), .Y(n5062) );
  MUX2X1 U5235 ( .B(n5066), .A(n5067), .S(n6242), .Y(n5065) );
  MUX2X1 U5236 ( .B(n5069), .A(n5070), .S(n6305), .Y(n5068) );
  MUX2X1 U5237 ( .B(n5072), .A(n5073), .S(n6306), .Y(n5071) );
  MUX2X1 U5238 ( .B(n5075), .A(n5076), .S(n6306), .Y(n5074) );
  MUX2X1 U5239 ( .B(n5078), .A(n5079), .S(n6306), .Y(n5077) );
  MUX2X1 U5240 ( .B(n5081), .A(n5082), .S(n6242), .Y(n5080) );
  MUX2X1 U5241 ( .B(n5084), .A(n5085), .S(n6306), .Y(n5083) );
  MUX2X1 U5242 ( .B(n5087), .A(n5088), .S(n6306), .Y(n5086) );
  MUX2X1 U5243 ( .B(n5090), .A(n5091), .S(n6306), .Y(n5089) );
  MUX2X1 U5244 ( .B(n5093), .A(n5094), .S(n6306), .Y(n5092) );
  MUX2X1 U5245 ( .B(n5096), .A(n5097), .S(n6242), .Y(n5095) );
  MUX2X1 U5246 ( .B(n5099), .A(n5100), .S(n6306), .Y(n5098) );
  MUX2X1 U5247 ( .B(n5102), .A(n5103), .S(n6306), .Y(n5101) );
  MUX2X1 U5248 ( .B(n5105), .A(n5106), .S(n6306), .Y(n5104) );
  MUX2X1 U5249 ( .B(n5108), .A(n5109), .S(n6306), .Y(n5107) );
  MUX2X1 U5250 ( .B(n5111), .A(n5112), .S(n6242), .Y(n5110) );
  MUX2X1 U5251 ( .B(n5113), .A(n5114), .S(n6232), .Y(N99) );
  MUX2X1 U5252 ( .B(n5116), .A(n5117), .S(n6306), .Y(n5115) );
  MUX2X1 U5253 ( .B(n5119), .A(n5120), .S(n6306), .Y(n5118) );
  MUX2X1 U5254 ( .B(n5122), .A(n5123), .S(n6307), .Y(n5121) );
  MUX2X1 U5255 ( .B(n5125), .A(n5126), .S(n6307), .Y(n5124) );
  MUX2X1 U5256 ( .B(n5128), .A(n5129), .S(n6242), .Y(n5127) );
  MUX2X1 U5257 ( .B(n5131), .A(n5132), .S(n6307), .Y(n5130) );
  MUX2X1 U5258 ( .B(n5134), .A(n5135), .S(n6307), .Y(n5133) );
  MUX2X1 U5259 ( .B(n5137), .A(n5138), .S(n6307), .Y(n5136) );
  MUX2X1 U5260 ( .B(n5140), .A(n5141), .S(n6307), .Y(n5139) );
  MUX2X1 U5261 ( .B(n5143), .A(n5144), .S(n6242), .Y(n5142) );
  MUX2X1 U5262 ( .B(n5146), .A(n5147), .S(n6307), .Y(n5145) );
  MUX2X1 U5263 ( .B(n5149), .A(n5150), .S(n6307), .Y(n5148) );
  MUX2X1 U5264 ( .B(n5152), .A(n5153), .S(n6307), .Y(n5151) );
  MUX2X1 U5265 ( .B(n5155), .A(n5156), .S(n6307), .Y(n5154) );
  MUX2X1 U5266 ( .B(n5158), .A(n5159), .S(n6242), .Y(n5157) );
  MUX2X1 U5267 ( .B(n5161), .A(n5162), .S(n6307), .Y(n5160) );
  MUX2X1 U5268 ( .B(n5164), .A(n5165), .S(n6307), .Y(n5163) );
  MUX2X1 U5269 ( .B(n5167), .A(n5168), .S(n6307), .Y(n5166) );
  MUX2X1 U5270 ( .B(n5170), .A(n5171), .S(n6308), .Y(n5169) );
  MUX2X1 U5271 ( .B(n5173), .A(n5174), .S(n6242), .Y(n5172) );
  MUX2X1 U5272 ( .B(n5175), .A(n5176), .S(n6232), .Y(N98) );
  MUX2X1 U5273 ( .B(n5178), .A(n5179), .S(n6308), .Y(n5177) );
  MUX2X1 U5274 ( .B(n5181), .A(n5182), .S(n6308), .Y(n5180) );
  MUX2X1 U5275 ( .B(n5184), .A(n5185), .S(n6308), .Y(n5183) );
  MUX2X1 U5276 ( .B(n5187), .A(n5188), .S(n6308), .Y(n5186) );
  MUX2X1 U5277 ( .B(n5190), .A(n5191), .S(n6242), .Y(n5189) );
  MUX2X1 U5278 ( .B(n5193), .A(n5194), .S(n6308), .Y(n5192) );
  MUX2X1 U5279 ( .B(n5196), .A(n5197), .S(n6308), .Y(n5195) );
  MUX2X1 U5280 ( .B(n5199), .A(n5200), .S(n6308), .Y(n5198) );
  MUX2X1 U5281 ( .B(n5202), .A(n5203), .S(n6308), .Y(n5201) );
  MUX2X1 U5282 ( .B(n5205), .A(n5206), .S(n6242), .Y(n5204) );
  MUX2X1 U5283 ( .B(n5208), .A(n5209), .S(n6308), .Y(n5207) );
  MUX2X1 U5284 ( .B(n5211), .A(n5212), .S(n6308), .Y(n5210) );
  MUX2X1 U5285 ( .B(n5214), .A(n5215), .S(n6308), .Y(n5213) );
  MUX2X1 U5286 ( .B(n5217), .A(n5218), .S(n6308), .Y(n5216) );
  MUX2X1 U5287 ( .B(n5220), .A(n5221), .S(n6242), .Y(n5219) );
  MUX2X1 U5288 ( .B(n5223), .A(n5224), .S(n6309), .Y(n5222) );
  MUX2X1 U5289 ( .B(n5226), .A(n5227), .S(n6309), .Y(n5225) );
  MUX2X1 U5290 ( .B(n5229), .A(n5230), .S(n6309), .Y(n5228) );
  MUX2X1 U5291 ( .B(n5232), .A(n5233), .S(n6309), .Y(n5231) );
  MUX2X1 U5292 ( .B(n5235), .A(n5236), .S(n6243), .Y(n5234) );
  MUX2X1 U5293 ( .B(n5237), .A(n5238), .S(n6232), .Y(N97) );
  MUX2X1 U5294 ( .B(n5240), .A(n5241), .S(n6309), .Y(n5239) );
  MUX2X1 U5295 ( .B(n5243), .A(n5244), .S(n6309), .Y(n5242) );
  MUX2X1 U5296 ( .B(n5246), .A(n5247), .S(n6309), .Y(n5245) );
  MUX2X1 U5297 ( .B(n5249), .A(n5250), .S(n6309), .Y(n5248) );
  MUX2X1 U5298 ( .B(n5252), .A(n5253), .S(n6243), .Y(n5251) );
  MUX2X1 U5299 ( .B(n5255), .A(n5256), .S(n6309), .Y(n5254) );
  MUX2X1 U5300 ( .B(n5258), .A(n5259), .S(n6309), .Y(n5257) );
  MUX2X1 U5301 ( .B(n5261), .A(n5262), .S(n6309), .Y(n5260) );
  MUX2X1 U5302 ( .B(n5264), .A(n5265), .S(n6309), .Y(n5263) );
  MUX2X1 U5303 ( .B(n5267), .A(n5268), .S(n6243), .Y(n5266) );
  MUX2X1 U5304 ( .B(n5270), .A(n5271), .S(n6309), .Y(n5269) );
  MUX2X1 U5305 ( .B(n5273), .A(n5274), .S(n6310), .Y(n5272) );
  MUX2X1 U5306 ( .B(n5276), .A(n5277), .S(n6310), .Y(n5275) );
  MUX2X1 U5307 ( .B(n5279), .A(n5280), .S(n6310), .Y(n5278) );
  MUX2X1 U5308 ( .B(n5282), .A(n5283), .S(n6243), .Y(n5281) );
  MUX2X1 U5309 ( .B(n5285), .A(n5286), .S(n6310), .Y(n5284) );
  MUX2X1 U5310 ( .B(n5288), .A(n5289), .S(n6310), .Y(n5287) );
  MUX2X1 U5311 ( .B(n5291), .A(n5292), .S(n6310), .Y(n5290) );
  MUX2X1 U5312 ( .B(n5294), .A(n5295), .S(n6310), .Y(n5293) );
  MUX2X1 U5313 ( .B(n5297), .A(n5298), .S(n6243), .Y(n5296) );
  MUX2X1 U5314 ( .B(n5299), .A(n5300), .S(n6232), .Y(N96) );
  MUX2X1 U5315 ( .B(n5302), .A(n5303), .S(n6310), .Y(n5301) );
  MUX2X1 U5316 ( .B(n5305), .A(n5306), .S(n6310), .Y(n5304) );
  MUX2X1 U5317 ( .B(n5308), .A(n5309), .S(n6310), .Y(n5307) );
  MUX2X1 U5318 ( .B(n5311), .A(n5312), .S(n6310), .Y(n5310) );
  MUX2X1 U5319 ( .B(n5314), .A(n5315), .S(n6243), .Y(n5313) );
  MUX2X1 U5320 ( .B(n5317), .A(n5318), .S(n6310), .Y(n5316) );
  MUX2X1 U5321 ( .B(n5320), .A(n5321), .S(n6310), .Y(n5319) );
  MUX2X1 U5322 ( .B(n5323), .A(n5324), .S(n6311), .Y(n5322) );
  MUX2X1 U5323 ( .B(n5326), .A(n5327), .S(n6311), .Y(n5325) );
  MUX2X1 U5324 ( .B(n5329), .A(n5330), .S(n6243), .Y(n5328) );
  MUX2X1 U5325 ( .B(n5332), .A(n5333), .S(n6311), .Y(n5331) );
  MUX2X1 U5326 ( .B(n5335), .A(n5336), .S(n6311), .Y(n5334) );
  MUX2X1 U5327 ( .B(n5338), .A(n5339), .S(n6311), .Y(n5337) );
  MUX2X1 U5328 ( .B(n5341), .A(n5342), .S(n6311), .Y(n5340) );
  MUX2X1 U5329 ( .B(n5344), .A(n5345), .S(n6243), .Y(n5343) );
  MUX2X1 U5330 ( .B(n5347), .A(n5348), .S(n6311), .Y(n5346) );
  MUX2X1 U5331 ( .B(n5350), .A(n5351), .S(n6311), .Y(n5349) );
  MUX2X1 U5332 ( .B(n5353), .A(n5354), .S(n6311), .Y(n5352) );
  MUX2X1 U5333 ( .B(n5356), .A(n5357), .S(n6311), .Y(n5355) );
  MUX2X1 U5334 ( .B(n5359), .A(n5360), .S(n6243), .Y(n5358) );
  MUX2X1 U5335 ( .B(n5361), .A(n5362), .S(n6232), .Y(N95) );
  MUX2X1 U5336 ( .B(n5364), .A(n5365), .S(n6311), .Y(n5363) );
  MUX2X1 U5337 ( .B(n5367), .A(n5368), .S(n6311), .Y(n5366) );
  MUX2X1 U5338 ( .B(n5370), .A(n5371), .S(n6311), .Y(n5369) );
  MUX2X1 U5339 ( .B(n5373), .A(n5374), .S(n6312), .Y(n5372) );
  MUX2X1 U5340 ( .B(n5376), .A(n5377), .S(n6243), .Y(n5375) );
  MUX2X1 U5341 ( .B(n5379), .A(n5380), .S(n6312), .Y(n5378) );
  MUX2X1 U5342 ( .B(n5382), .A(n5383), .S(n6312), .Y(n5381) );
  MUX2X1 U5343 ( .B(n5385), .A(n5386), .S(n6312), .Y(n5384) );
  MUX2X1 U5344 ( .B(n5388), .A(n5389), .S(n6312), .Y(n5387) );
  MUX2X1 U5345 ( .B(n5391), .A(n5392), .S(n6243), .Y(n5390) );
  MUX2X1 U5346 ( .B(n5394), .A(n5395), .S(n6312), .Y(n5393) );
  MUX2X1 U5347 ( .B(n5397), .A(n5398), .S(n6312), .Y(n5396) );
  MUX2X1 U5348 ( .B(n5400), .A(n5401), .S(n6312), .Y(n5399) );
  MUX2X1 U5349 ( .B(n5403), .A(n5404), .S(n6312), .Y(n5402) );
  MUX2X1 U5350 ( .B(n5406), .A(n5407), .S(n6243), .Y(n5405) );
  MUX2X1 U5351 ( .B(n5409), .A(n5410), .S(n6312), .Y(n5408) );
  MUX2X1 U5352 ( .B(n5412), .A(n5413), .S(n6312), .Y(n5411) );
  MUX2X1 U5353 ( .B(n5415), .A(n5416), .S(n6312), .Y(n5414) );
  MUX2X1 U5354 ( .B(n5418), .A(n5419), .S(n6312), .Y(n5417) );
  MUX2X1 U5355 ( .B(n5421), .A(n5422), .S(n6243), .Y(n5420) );
  MUX2X1 U5356 ( .B(n5423), .A(n5424), .S(n6232), .Y(N94) );
  MUX2X1 U5357 ( .B(n5426), .A(n5427), .S(n6313), .Y(n5425) );
  MUX2X1 U5358 ( .B(n5429), .A(n5430), .S(n6313), .Y(n5428) );
  MUX2X1 U5359 ( .B(n5432), .A(n5433), .S(n6313), .Y(n5431) );
  MUX2X1 U5360 ( .B(n5435), .A(n5436), .S(n6313), .Y(n5434) );
  MUX2X1 U5361 ( .B(n5438), .A(n5439), .S(n6244), .Y(n5437) );
  MUX2X1 U5362 ( .B(n5441), .A(n5442), .S(n6313), .Y(n5440) );
  MUX2X1 U5363 ( .B(n5444), .A(n5445), .S(n6313), .Y(n5443) );
  MUX2X1 U5364 ( .B(n5447), .A(n5448), .S(n6313), .Y(n5446) );
  MUX2X1 U5365 ( .B(n5450), .A(n5451), .S(n6313), .Y(n5449) );
  MUX2X1 U5366 ( .B(n5453), .A(n5454), .S(n6244), .Y(n5452) );
  MUX2X1 U5367 ( .B(n5456), .A(n5457), .S(n6313), .Y(n5455) );
  MUX2X1 U5368 ( .B(n5459), .A(n5460), .S(n6313), .Y(n5458) );
  MUX2X1 U5369 ( .B(n5462), .A(n5463), .S(n6313), .Y(n5461) );
  MUX2X1 U5370 ( .B(n5465), .A(n5466), .S(n6313), .Y(n5464) );
  MUX2X1 U5371 ( .B(n5468), .A(n5469), .S(n6244), .Y(n5467) );
  MUX2X1 U5372 ( .B(n5471), .A(n5472), .S(n6313), .Y(n5470) );
  MUX2X1 U5373 ( .B(n5474), .A(n5475), .S(n6314), .Y(n5473) );
  MUX2X1 U5374 ( .B(n5477), .A(n5478), .S(n6314), .Y(n5476) );
  MUX2X1 U5375 ( .B(n5480), .A(n5481), .S(n6314), .Y(n5479) );
  MUX2X1 U5376 ( .B(n5483), .A(n5484), .S(n6244), .Y(n5482) );
  MUX2X1 U5377 ( .B(n5485), .A(n5486), .S(N15), .Y(N93) );
  MUX2X1 U5378 ( .B(n5488), .A(n5489), .S(n6314), .Y(n5487) );
  MUX2X1 U5379 ( .B(n5491), .A(n5492), .S(n6314), .Y(n5490) );
  MUX2X1 U5380 ( .B(n5494), .A(n5495), .S(n6314), .Y(n5493) );
  MUX2X1 U5381 ( .B(n5497), .A(n5498), .S(n6314), .Y(n5496) );
  MUX2X1 U5382 ( .B(n5500), .A(n5501), .S(n6244), .Y(n5499) );
  MUX2X1 U5383 ( .B(n5503), .A(n5504), .S(n6314), .Y(n5502) );
  MUX2X1 U5384 ( .B(n5506), .A(n5507), .S(n6314), .Y(n5505) );
  MUX2X1 U5385 ( .B(n5509), .A(n5510), .S(n6314), .Y(n5508) );
  MUX2X1 U5386 ( .B(n5512), .A(n5513), .S(n6314), .Y(n5511) );
  MUX2X1 U5387 ( .B(n5515), .A(n5516), .S(n6244), .Y(n5514) );
  MUX2X1 U5388 ( .B(n5518), .A(n5519), .S(n6314), .Y(n5517) );
  MUX2X1 U5389 ( .B(n5521), .A(n5522), .S(n6314), .Y(n5520) );
  MUX2X1 U5390 ( .B(n5524), .A(n5525), .S(n6315), .Y(n5523) );
  MUX2X1 U5391 ( .B(n5527), .A(n5528), .S(n6315), .Y(n5526) );
  MUX2X1 U5392 ( .B(n5530), .A(n5531), .S(n6244), .Y(n5529) );
  MUX2X1 U5393 ( .B(n5533), .A(n5534), .S(n6315), .Y(n5532) );
  MUX2X1 U5394 ( .B(n5536), .A(n5537), .S(n6315), .Y(n5535) );
  MUX2X1 U5395 ( .B(n5539), .A(n5540), .S(n6315), .Y(n5538) );
  MUX2X1 U5396 ( .B(n5542), .A(n5543), .S(n6315), .Y(n5541) );
  MUX2X1 U5397 ( .B(n5545), .A(n5546), .S(n6244), .Y(n5544) );
  MUX2X1 U5398 ( .B(n5547), .A(n5548), .S(N15), .Y(N92) );
  MUX2X1 U5399 ( .B(n5550), .A(n5551), .S(n6315), .Y(n5549) );
  MUX2X1 U5400 ( .B(n5553), .A(n5554), .S(n6315), .Y(n5552) );
  MUX2X1 U5401 ( .B(n5556), .A(n5557), .S(n6315), .Y(n5555) );
  MUX2X1 U5402 ( .B(n5559), .A(n5560), .S(n6315), .Y(n5558) );
  MUX2X1 U5403 ( .B(n5562), .A(n5563), .S(n6244), .Y(n5561) );
  MUX2X1 U5404 ( .B(n5565), .A(n5566), .S(n6315), .Y(n5564) );
  MUX2X1 U5405 ( .B(n5568), .A(n5569), .S(n6315), .Y(n5567) );
  MUX2X1 U5406 ( .B(n5571), .A(n5572), .S(n6315), .Y(n5570) );
  MUX2X1 U5407 ( .B(n5574), .A(n5575), .S(n6316), .Y(n5573) );
  MUX2X1 U5408 ( .B(n5577), .A(n5578), .S(n6244), .Y(n5576) );
  MUX2X1 U5409 ( .B(n5580), .A(n5581), .S(n6316), .Y(n5579) );
  MUX2X1 U5410 ( .B(n5583), .A(n5584), .S(n6316), .Y(n5582) );
  MUX2X1 U5411 ( .B(n5586), .A(n5587), .S(n6316), .Y(n5585) );
  MUX2X1 U5412 ( .B(n5589), .A(n5590), .S(n6316), .Y(n5588) );
  MUX2X1 U5413 ( .B(n5592), .A(n5593), .S(n6244), .Y(n5591) );
  MUX2X1 U5414 ( .B(n5595), .A(n5596), .S(n6316), .Y(n5594) );
  MUX2X1 U5415 ( .B(n5598), .A(n5599), .S(n6316), .Y(n5597) );
  MUX2X1 U5416 ( .B(n5601), .A(n5602), .S(n6316), .Y(n5600) );
  MUX2X1 U5417 ( .B(n5604), .A(n5605), .S(n6316), .Y(n5603) );
  MUX2X1 U5418 ( .B(n5607), .A(n5608), .S(n6244), .Y(n5606) );
  MUX2X1 U5419 ( .B(n5609), .A(n5610), .S(N15), .Y(N91) );
  MUX2X1 U5420 ( .B(n5612), .A(n5613), .S(n6316), .Y(n5611) );
  MUX2X1 U5421 ( .B(n5615), .A(n5616), .S(n6316), .Y(n5614) );
  MUX2X1 U5422 ( .B(n5618), .A(n5619), .S(n6316), .Y(n5617) );
  MUX2X1 U5423 ( .B(n5621), .A(n5622), .S(n6316), .Y(n5620) );
  MUX2X1 U5424 ( .B(n5624), .A(n5625), .S(n6244), .Y(n5623) );
  MUX2X1 U5425 ( .B(n5627), .A(n5628), .S(n6317), .Y(n5626) );
  MUX2X1 U5426 ( .B(n5630), .A(n5631), .S(n6317), .Y(n5629) );
  MUX2X1 U5427 ( .B(n5633), .A(n5634), .S(n6317), .Y(n5632) );
  MUX2X1 U5428 ( .B(n5636), .A(n5637), .S(n6317), .Y(n5635) );
  MUX2X1 U5429 ( .B(n5639), .A(n5640), .S(n6245), .Y(n5638) );
  MUX2X1 U5430 ( .B(n5642), .A(n5643), .S(n6317), .Y(n5641) );
  MUX2X1 U5431 ( .B(n5645), .A(n5646), .S(n6317), .Y(n5644) );
  MUX2X1 U5432 ( .B(n5648), .A(n5649), .S(n6317), .Y(n5647) );
  MUX2X1 U5433 ( .B(n5651), .A(n5652), .S(n6317), .Y(n5650) );
  MUX2X1 U5434 ( .B(n5654), .A(n5655), .S(n6245), .Y(n5653) );
  MUX2X1 U5435 ( .B(n5657), .A(n5658), .S(n6317), .Y(n5656) );
  MUX2X1 U5436 ( .B(n5660), .A(n5661), .S(n6317), .Y(n5659) );
  MUX2X1 U5437 ( .B(n5663), .A(n5664), .S(n6317), .Y(n5662) );
  MUX2X1 U5438 ( .B(n5666), .A(n5667), .S(n6317), .Y(n5665) );
  MUX2X1 U5439 ( .B(n5669), .A(n5670), .S(n6245), .Y(n5668) );
  MUX2X1 U5440 ( .B(n5671), .A(n5672), .S(n6232), .Y(N90) );
  MUX2X1 U5441 ( .B(n5674), .A(n5675), .S(n6317), .Y(n5673) );
  MUX2X1 U5442 ( .B(n5677), .A(n5678), .S(n6318), .Y(n5676) );
  MUX2X1 U5443 ( .B(n5680), .A(n5681), .S(n6318), .Y(n5679) );
  MUX2X1 U5444 ( .B(n5683), .A(n5684), .S(n6318), .Y(n5682) );
  MUX2X1 U5445 ( .B(n5686), .A(n5687), .S(n6245), .Y(n5685) );
  MUX2X1 U5446 ( .B(n5689), .A(n5690), .S(n6318), .Y(n5688) );
  MUX2X1 U5447 ( .B(n5692), .A(n5693), .S(n6318), .Y(n5691) );
  MUX2X1 U5448 ( .B(n5695), .A(n5696), .S(n6318), .Y(n5694) );
  MUX2X1 U5449 ( .B(n5698), .A(n5699), .S(n6318), .Y(n5697) );
  MUX2X1 U5450 ( .B(n5701), .A(n5702), .S(n6245), .Y(n5700) );
  MUX2X1 U5451 ( .B(n5704), .A(n5705), .S(n6318), .Y(n5703) );
  MUX2X1 U5452 ( .B(n5707), .A(n5708), .S(n6318), .Y(n5706) );
  MUX2X1 U5453 ( .B(n5710), .A(n5711), .S(n6318), .Y(n5709) );
  MUX2X1 U5454 ( .B(n5713), .A(n5714), .S(n6318), .Y(n5712) );
  MUX2X1 U5455 ( .B(n5716), .A(n5717), .S(n6245), .Y(n5715) );
  MUX2X1 U5456 ( .B(n5719), .A(n5720), .S(n6318), .Y(n5718) );
  MUX2X1 U5457 ( .B(n5722), .A(n5723), .S(n6318), .Y(n5721) );
  MUX2X1 U5458 ( .B(n5725), .A(n5726), .S(n6319), .Y(n5724) );
  MUX2X1 U5459 ( .B(n5728), .A(n5729), .S(n6319), .Y(n5727) );
  MUX2X1 U5460 ( .B(n5731), .A(n5732), .S(n6245), .Y(n5730) );
  MUX2X1 U5461 ( .B(n5733), .A(n5734), .S(n6232), .Y(N89) );
  MUX2X1 U5462 ( .B(n5736), .A(n5737), .S(n6319), .Y(n5735) );
  MUX2X1 U5463 ( .B(n5739), .A(n5740), .S(n6319), .Y(n5738) );
  MUX2X1 U5464 ( .B(n5742), .A(n5743), .S(n6319), .Y(n5741) );
  MUX2X1 U5465 ( .B(n5745), .A(n5746), .S(n6319), .Y(n5744) );
  MUX2X1 U5466 ( .B(n5748), .A(n5749), .S(n6245), .Y(n5747) );
  MUX2X1 U5467 ( .B(n5751), .A(n5752), .S(n6319), .Y(n5750) );
  MUX2X1 U5468 ( .B(n5754), .A(n5755), .S(n6319), .Y(n5753) );
  MUX2X1 U5469 ( .B(n5757), .A(n5758), .S(n6319), .Y(n5756) );
  MUX2X1 U5470 ( .B(n5760), .A(n5761), .S(n6319), .Y(n5759) );
  MUX2X1 U5471 ( .B(n5763), .A(n5764), .S(n6245), .Y(n5762) );
  MUX2X1 U5472 ( .B(n5766), .A(n5767), .S(n6319), .Y(n5765) );
  MUX2X1 U5473 ( .B(n5769), .A(n5770), .S(n6319), .Y(n5768) );
  MUX2X1 U5474 ( .B(n5772), .A(n5773), .S(n6319), .Y(n5771) );
  MUX2X1 U5475 ( .B(n5775), .A(n5776), .S(n6320), .Y(n5774) );
  MUX2X1 U5476 ( .B(n5778), .A(n5779), .S(n6245), .Y(n5777) );
  MUX2X1 U5477 ( .B(n5781), .A(n5782), .S(n6320), .Y(n5780) );
  MUX2X1 U5478 ( .B(n5784), .A(n5785), .S(n6320), .Y(n5783) );
  MUX2X1 U5479 ( .B(n5787), .A(n5788), .S(n6320), .Y(n5786) );
  MUX2X1 U5480 ( .B(n5790), .A(n5791), .S(n6320), .Y(n5789) );
  MUX2X1 U5481 ( .B(n5793), .A(n5794), .S(n6245), .Y(n5792) );
  MUX2X1 U5482 ( .B(n5795), .A(n5796), .S(n6232), .Y(N88) );
  MUX2X1 U5483 ( .B(n5798), .A(n5799), .S(n6320), .Y(n5797) );
  MUX2X1 U5484 ( .B(n5801), .A(n5802), .S(n6320), .Y(n5800) );
  MUX2X1 U5485 ( .B(n5804), .A(n5805), .S(n6320), .Y(n5803) );
  MUX2X1 U5486 ( .B(n5807), .A(n5808), .S(n6320), .Y(n5806) );
  MUX2X1 U5487 ( .B(n5810), .A(n5811), .S(n6245), .Y(n5809) );
  MUX2X1 U5488 ( .B(n5813), .A(n5814), .S(n6320), .Y(n5812) );
  MUX2X1 U5489 ( .B(n5816), .A(n5817), .S(n6320), .Y(n5815) );
  MUX2X1 U5490 ( .B(n5819), .A(n5820), .S(n6320), .Y(n5818) );
  MUX2X1 U5491 ( .B(n5822), .A(n5823), .S(n6320), .Y(n5821) );
  MUX2X1 U5492 ( .B(n5825), .A(n5826), .S(n6245), .Y(n5824) );
  MUX2X1 U5493 ( .B(n5828), .A(n5829), .S(n6321), .Y(n5827) );
  MUX2X1 U5494 ( .B(n5831), .A(n5832), .S(n6321), .Y(n5830) );
  MUX2X1 U5495 ( .B(n5834), .A(n5835), .S(n6321), .Y(n5833) );
  MUX2X1 U5496 ( .B(n5837), .A(n5838), .S(n6321), .Y(n5836) );
  MUX2X1 U5497 ( .B(n5840), .A(n5841), .S(n6246), .Y(n5839) );
  MUX2X1 U5498 ( .B(n5843), .A(n5844), .S(n6321), .Y(n5842) );
  MUX2X1 U5499 ( .B(n5846), .A(n5847), .S(n6321), .Y(n5845) );
  MUX2X1 U5500 ( .B(n5849), .A(n5850), .S(n6321), .Y(n5848) );
  MUX2X1 U5501 ( .B(n5852), .A(n5853), .S(n6321), .Y(n5851) );
  MUX2X1 U5502 ( .B(n5855), .A(n5856), .S(n6246), .Y(n5854) );
  MUX2X1 U5503 ( .B(n5857), .A(n5858), .S(n6232), .Y(N87) );
  MUX2X1 U5504 ( .B(n5860), .A(n5861), .S(n6321), .Y(n5859) );
  MUX2X1 U5505 ( .B(n5863), .A(n5864), .S(n6321), .Y(n5862) );
  MUX2X1 U5506 ( .B(n5866), .A(n5867), .S(n6321), .Y(n5865) );
  MUX2X1 U5507 ( .B(n5869), .A(n5870), .S(n6321), .Y(n5868) );
  MUX2X1 U5508 ( .B(n5872), .A(n5873), .S(n6246), .Y(n5871) );
  MUX2X1 U5509 ( .B(n5875), .A(n5876), .S(n6321), .Y(n5874) );
  MUX2X1 U5510 ( .B(n5878), .A(n5879), .S(n6322), .Y(n5877) );
  MUX2X1 U5511 ( .B(n5881), .A(n5882), .S(n6322), .Y(n5880) );
  MUX2X1 U5512 ( .B(n5884), .A(n5885), .S(n6322), .Y(n5883) );
  MUX2X1 U5513 ( .B(n5887), .A(n5888), .S(n6246), .Y(n5886) );
  MUX2X1 U5514 ( .B(n5890), .A(n5891), .S(n6322), .Y(n5889) );
  MUX2X1 U5515 ( .B(n5893), .A(n5894), .S(n6322), .Y(n5892) );
  MUX2X1 U5516 ( .B(n5896), .A(n5897), .S(n6322), .Y(n5895) );
  MUX2X1 U5517 ( .B(n5899), .A(n5900), .S(n6322), .Y(n5898) );
  MUX2X1 U5518 ( .B(n5902), .A(n5903), .S(n6246), .Y(n5901) );
  MUX2X1 U5519 ( .B(n5905), .A(n5906), .S(n6322), .Y(n5904) );
  MUX2X1 U5520 ( .B(n5908), .A(n5909), .S(n6322), .Y(n5907) );
  MUX2X1 U5521 ( .B(n5911), .A(n5912), .S(n6322), .Y(n5910) );
  MUX2X1 U5522 ( .B(n5914), .A(n5915), .S(n6322), .Y(n5913) );
  MUX2X1 U5523 ( .B(n5917), .A(n5918), .S(n6246), .Y(n5916) );
  MUX2X1 U5524 ( .B(n5919), .A(n5920), .S(n6232), .Y(N86) );
  MUX2X1 U5525 ( .B(n5922), .A(n5923), .S(n6322), .Y(n5921) );
  MUX2X1 U5526 ( .B(n5925), .A(n5926), .S(n6322), .Y(n5924) );
  MUX2X1 U5527 ( .B(n5928), .A(n5929), .S(n6323), .Y(n5927) );
  MUX2X1 U5528 ( .B(n5931), .A(n5932), .S(n6323), .Y(n5930) );
  MUX2X1 U5529 ( .B(n5934), .A(n5935), .S(n6246), .Y(n5933) );
  MUX2X1 U5530 ( .B(n5937), .A(n5938), .S(n6323), .Y(n5936) );
  MUX2X1 U5531 ( .B(n5940), .A(n5941), .S(n6323), .Y(n5939) );
  MUX2X1 U5532 ( .B(n5943), .A(n5944), .S(n6323), .Y(n5942) );
  MUX2X1 U5533 ( .B(n5946), .A(n5947), .S(n6323), .Y(n5945) );
  MUX2X1 U5534 ( .B(n5949), .A(n5950), .S(n6246), .Y(n5948) );
  MUX2X1 U5535 ( .B(n5952), .A(n5953), .S(n6323), .Y(n5951) );
  MUX2X1 U5536 ( .B(n5955), .A(n5956), .S(n6323), .Y(n5954) );
  MUX2X1 U5537 ( .B(n5958), .A(n5959), .S(n6323), .Y(n5957) );
  MUX2X1 U5538 ( .B(n5961), .A(n5962), .S(n6323), .Y(n5960) );
  MUX2X1 U5539 ( .B(n5964), .A(n5965), .S(n6246), .Y(n5963) );
  MUX2X1 U5540 ( .B(n5967), .A(n5968), .S(n6323), .Y(n5966) );
  MUX2X1 U5541 ( .B(n5970), .A(n5971), .S(n6323), .Y(n5969) );
  MUX2X1 U5542 ( .B(n5973), .A(n5974), .S(n6323), .Y(n5972) );
  MUX2X1 U5543 ( .B(n5976), .A(n5977), .S(n6324), .Y(n5975) );
  MUX2X1 U5544 ( .B(n5979), .A(n5980), .S(n6246), .Y(n5978) );
  MUX2X1 U5545 ( .B(n5981), .A(n5982), .S(n6232), .Y(N85) );
  MUX2X1 U5546 ( .B(n5984), .A(n5985), .S(n6324), .Y(n5983) );
  MUX2X1 U5547 ( .B(n5987), .A(n5988), .S(n6324), .Y(n5986) );
  MUX2X1 U5548 ( .B(n5990), .A(n5991), .S(n6324), .Y(n5989) );
  MUX2X1 U5549 ( .B(n5993), .A(n5994), .S(n6324), .Y(n5992) );
  MUX2X1 U5550 ( .B(n5996), .A(n5997), .S(n6246), .Y(n5995) );
  MUX2X1 U5551 ( .B(n5999), .A(n6000), .S(n6324), .Y(n5998) );
  MUX2X1 U5552 ( .B(n6002), .A(n6003), .S(n6324), .Y(n6001) );
  MUX2X1 U5553 ( .B(n6005), .A(n6006), .S(n6324), .Y(n6004) );
  MUX2X1 U5554 ( .B(n6008), .A(n6009), .S(n6324), .Y(n6007) );
  MUX2X1 U5555 ( .B(n6011), .A(n6012), .S(n6246), .Y(n6010) );
  MUX2X1 U5556 ( .B(n6014), .A(n6015), .S(n6324), .Y(n6013) );
  MUX2X1 U5557 ( .B(n6017), .A(n6018), .S(n6324), .Y(n6016) );
  MUX2X1 U5558 ( .B(n6020), .A(n6021), .S(n6324), .Y(n6019) );
  MUX2X1 U5559 ( .B(n6023), .A(n6024), .S(n6324), .Y(n6022) );
  MUX2X1 U5560 ( .B(n6026), .A(n6027), .S(n6246), .Y(n6025) );
  MUX2X1 U5561 ( .B(n6029), .A(n6030), .S(n6325), .Y(n6028) );
  MUX2X1 U5562 ( .B(n6032), .A(n6033), .S(n6325), .Y(n6031) );
  MUX2X1 U5563 ( .B(n6035), .A(n6036), .S(n6325), .Y(n6034) );
  MUX2X1 U5564 ( .B(n6038), .A(n6039), .S(n6325), .Y(n6037) );
  MUX2X1 U5565 ( .B(n6041), .A(n6042), .S(n6247), .Y(n6040) );
  MUX2X1 U5566 ( .B(n6043), .A(n6044), .S(n6232), .Y(N84) );
  MUX2X1 U5567 ( .B(n6046), .A(n6047), .S(n6325), .Y(n6045) );
  MUX2X1 U5568 ( .B(n6049), .A(n6050), .S(n6325), .Y(n6048) );
  MUX2X1 U5569 ( .B(n6052), .A(n6053), .S(n6325), .Y(n6051) );
  MUX2X1 U5570 ( .B(n6055), .A(n6056), .S(n6325), .Y(n6054) );
  MUX2X1 U5571 ( .B(n6058), .A(n6059), .S(n6247), .Y(n6057) );
  MUX2X1 U5572 ( .B(n6061), .A(n6062), .S(n6325), .Y(n6060) );
  MUX2X1 U5573 ( .B(n6064), .A(n6065), .S(n6325), .Y(n6063) );
  MUX2X1 U5574 ( .B(n6067), .A(n6068), .S(n6325), .Y(n6066) );
  MUX2X1 U5575 ( .B(n6070), .A(n6071), .S(n6325), .Y(n6069) );
  MUX2X1 U5576 ( .B(n6073), .A(n6074), .S(n6247), .Y(n6072) );
  MUX2X1 U5577 ( .B(n6076), .A(n6077), .S(n6325), .Y(n6075) );
  MUX2X1 U5578 ( .B(n6079), .A(n6080), .S(n6326), .Y(n6078) );
  MUX2X1 U5579 ( .B(n6082), .A(n6083), .S(n6326), .Y(n6081) );
  MUX2X1 U5580 ( .B(n6085), .A(n6086), .S(n6326), .Y(n6084) );
  MUX2X1 U5581 ( .B(n6088), .A(n6089), .S(n6247), .Y(n6087) );
  MUX2X1 U5582 ( .B(n6091), .A(n6092), .S(n6326), .Y(n6090) );
  MUX2X1 U5583 ( .B(n6094), .A(n6095), .S(n6326), .Y(n6093) );
  MUX2X1 U5584 ( .B(n6097), .A(n6098), .S(n6326), .Y(n6096) );
  MUX2X1 U5585 ( .B(n6100), .A(n6101), .S(n6326), .Y(n6099) );
  MUX2X1 U5586 ( .B(n6103), .A(n6104), .S(n6247), .Y(n6102) );
  MUX2X1 U5587 ( .B(n6105), .A(n6106), .S(n6232), .Y(N83) );
  MUX2X1 U5588 ( .B(n6108), .A(n6109), .S(n6326), .Y(n6107) );
  MUX2X1 U5589 ( .B(n6111), .A(n6112), .S(n6326), .Y(n6110) );
  MUX2X1 U5590 ( .B(n6114), .A(n6115), .S(n6326), .Y(n6113) );
  MUX2X1 U5591 ( .B(n6117), .A(n6118), .S(n6326), .Y(n6116) );
  MUX2X1 U5592 ( .B(n6120), .A(n6121), .S(n6247), .Y(n6119) );
  MUX2X1 U5593 ( .B(n6123), .A(n6124), .S(n6326), .Y(n6122) );
  MUX2X1 U5594 ( .B(n6126), .A(n6127), .S(n6326), .Y(n6125) );
  MUX2X1 U5595 ( .B(n6129), .A(n6130), .S(n6327), .Y(n6128) );
  MUX2X1 U5596 ( .B(n6132), .A(n6133), .S(n6327), .Y(n6131) );
  MUX2X1 U5597 ( .B(n6135), .A(n6136), .S(n6247), .Y(n6134) );
  MUX2X1 U5598 ( .B(n6138), .A(n6139), .S(n6327), .Y(n6137) );
  MUX2X1 U5599 ( .B(n6141), .A(n6142), .S(n6327), .Y(n6140) );
  MUX2X1 U5600 ( .B(n6144), .A(n6145), .S(n6327), .Y(n6143) );
  MUX2X1 U5601 ( .B(n6147), .A(n6148), .S(n6327), .Y(n6146) );
  MUX2X1 U5602 ( .B(n6150), .A(n6151), .S(n6247), .Y(n6149) );
  MUX2X1 U5603 ( .B(n6153), .A(n6154), .S(n6327), .Y(n6152) );
  MUX2X1 U5604 ( .B(n6156), .A(n6157), .S(n6327), .Y(n6155) );
  MUX2X1 U5605 ( .B(n6159), .A(n6160), .S(n6327), .Y(n6158) );
  MUX2X1 U5606 ( .B(n6162), .A(n6163), .S(n6327), .Y(n6161) );
  MUX2X1 U5607 ( .B(n6165), .A(n6166), .S(n6247), .Y(n6164) );
  MUX2X1 U5608 ( .B(n6167), .A(n6168), .S(n6232), .Y(N82) );
  MUX2X1 U5609 ( .B(n6170), .A(n6171), .S(n6327), .Y(n6169) );
  MUX2X1 U5610 ( .B(n6173), .A(n6174), .S(n6327), .Y(n6172) );
  MUX2X1 U5611 ( .B(n6176), .A(n6177), .S(n6327), .Y(n6175) );
  MUX2X1 U5612 ( .B(n6179), .A(n6180), .S(n6328), .Y(n6178) );
  MUX2X1 U5613 ( .B(n6182), .A(n6183), .S(n6247), .Y(n6181) );
  MUX2X1 U5614 ( .B(n6185), .A(n6186), .S(n6328), .Y(n6184) );
  MUX2X1 U5615 ( .B(n6188), .A(n6189), .S(n6328), .Y(n6187) );
  MUX2X1 U5616 ( .B(n6191), .A(n6192), .S(n6328), .Y(n6190) );
  MUX2X1 U5617 ( .B(n6194), .A(n6195), .S(n6328), .Y(n6193) );
  MUX2X1 U5618 ( .B(n6197), .A(n6198), .S(n6247), .Y(n6196) );
  MUX2X1 U5619 ( .B(n6200), .A(n6201), .S(n6328), .Y(n6199) );
  MUX2X1 U5620 ( .B(n6203), .A(n6204), .S(n6328), .Y(n6202) );
  MUX2X1 U5621 ( .B(n6206), .A(n6207), .S(n6328), .Y(n6205) );
  MUX2X1 U5622 ( .B(n6209), .A(n6210), .S(n6328), .Y(n6208) );
  MUX2X1 U5623 ( .B(n6212), .A(n6213), .S(n6247), .Y(n6211) );
  MUX2X1 U5624 ( .B(n6215), .A(n6216), .S(n6328), .Y(n6214) );
  MUX2X1 U5625 ( .B(n6218), .A(n6219), .S(n6328), .Y(n6217) );
  MUX2X1 U5626 ( .B(n6221), .A(n6222), .S(n6328), .Y(n6220) );
  MUX2X1 U5627 ( .B(n6224), .A(n6225), .S(n6328), .Y(n6223) );
  MUX2X1 U5628 ( .B(n6227), .A(n6228), .S(n6247), .Y(n6226) );
  MUX2X1 U5629 ( .B(n6229), .A(n6230), .S(n6232), .Y(N81) );
  MUX2X1 U5630 ( .B(\Mem[62][0] ), .A(\Mem[63][0] ), .S(n6361), .Y(n150) );
  MUX2X1 U5631 ( .B(\Mem[60][0] ), .A(\Mem[61][0] ), .S(n6361), .Y(n116) );
  MUX2X1 U5632 ( .B(\Mem[58][0] ), .A(\Mem[59][0] ), .S(n6361), .Y(n252) );
  MUX2X1 U5633 ( .B(\Mem[56][0] ), .A(\Mem[57][0] ), .S(n6361), .Y(n218) );
  MUX2X1 U5634 ( .B(n184), .A(n115), .S(n6248), .Y(n1456) );
  MUX2X1 U5635 ( .B(\Mem[54][0] ), .A(\Mem[55][0] ), .S(n6361), .Y(n356) );
  MUX2X1 U5636 ( .B(\Mem[52][0] ), .A(\Mem[53][0] ), .S(n6361), .Y(n320) );
  MUX2X1 U5637 ( .B(\Mem[50][0] ), .A(\Mem[51][0] ), .S(n6361), .Y(n657) );
  MUX2X1 U5638 ( .B(\Mem[48][0] ), .A(\Mem[49][0] ), .S(n6361), .Y(n623) );
  MUX2X1 U5639 ( .B(n390), .A(n286), .S(n6248), .Y(n1190) );
  MUX2X1 U5640 ( .B(\Mem[46][0] ), .A(\Mem[47][0] ), .S(n6361), .Y(n1959) );
  MUX2X1 U5641 ( .B(\Mem[44][0] ), .A(\Mem[45][0] ), .S(n6361), .Y(n1956) );
  MUX2X1 U5642 ( .B(\Mem[42][0] ), .A(\Mem[43][0] ), .S(n6362), .Y(n2027) );
  MUX2X1 U5643 ( .B(\Mem[40][0] ), .A(\Mem[41][0] ), .S(n6362), .Y(n2026) );
  MUX2X1 U5644 ( .B(n2025), .A(n1722), .S(n6248), .Y(n2228) );
  MUX2X1 U5645 ( .B(\Mem[38][0] ), .A(\Mem[39][0] ), .S(n6362), .Y(n2222) );
  MUX2X1 U5646 ( .B(\Mem[36][0] ), .A(\Mem[37][0] ), .S(n6362), .Y(n2221) );
  MUX2X1 U5647 ( .B(\Mem[34][0] ), .A(\Mem[35][0] ), .S(n6362), .Y(n2225) );
  MUX2X1 U5648 ( .B(\Mem[32][0] ), .A(\Mem[33][0] ), .S(n6362), .Y(n2224) );
  MUX2X1 U5649 ( .B(n2223), .A(n2218), .S(n6248), .Y(n2227) );
  MUX2X1 U5650 ( .B(n2226), .A(n923), .S(n6233), .Y(n2260) );
  MUX2X1 U5651 ( .B(\Mem[30][0] ), .A(\Mem[31][0] ), .S(n6362), .Y(n2231) );
  MUX2X1 U5652 ( .B(\Mem[28][0] ), .A(\Mem[29][0] ), .S(n6362), .Y(n2230) );
  MUX2X1 U5653 ( .B(\Mem[26][0] ), .A(\Mem[27][0] ), .S(n6362), .Y(n2234) );
  MUX2X1 U5654 ( .B(\Mem[24][0] ), .A(\Mem[25][0] ), .S(n6362), .Y(n2233) );
  MUX2X1 U5655 ( .B(n2232), .A(n2229), .S(n6248), .Y(n2243) );
  MUX2X1 U5656 ( .B(\Mem[22][0] ), .A(\Mem[23][0] ), .S(n6362), .Y(n2237) );
  MUX2X1 U5657 ( .B(\Mem[20][0] ), .A(\Mem[21][0] ), .S(n6362), .Y(n2236) );
  MUX2X1 U5658 ( .B(\Mem[18][0] ), .A(\Mem[19][0] ), .S(n6362), .Y(n2240) );
  MUX2X1 U5659 ( .B(\Mem[16][0] ), .A(\Mem[17][0] ), .S(n6363), .Y(n2239) );
  MUX2X1 U5660 ( .B(n2238), .A(n2235), .S(n6248), .Y(n2242) );
  MUX2X1 U5661 ( .B(\Mem[14][0] ), .A(\Mem[15][0] ), .S(n6363), .Y(n2246) );
  MUX2X1 U5662 ( .B(\Mem[12][0] ), .A(\Mem[13][0] ), .S(n6363), .Y(n2245) );
  MUX2X1 U5663 ( .B(\Mem[10][0] ), .A(\Mem[11][0] ), .S(n6363), .Y(n2249) );
  MUX2X1 U5664 ( .B(\Mem[8][0] ), .A(\Mem[9][0] ), .S(n6363), .Y(n2248) );
  MUX2X1 U5665 ( .B(n2247), .A(n2244), .S(n6248), .Y(n2258) );
  MUX2X1 U5666 ( .B(\Mem[6][0] ), .A(\Mem[7][0] ), .S(n6363), .Y(n2252) );
  MUX2X1 U5667 ( .B(\Mem[4][0] ), .A(\Mem[5][0] ), .S(n6363), .Y(n2251) );
  MUX2X1 U5668 ( .B(\Mem[2][0] ), .A(\Mem[3][0] ), .S(n6363), .Y(n2255) );
  MUX2X1 U5669 ( .B(\Mem[0][0] ), .A(\Mem[1][0] ), .S(n6363), .Y(n2254) );
  MUX2X1 U5670 ( .B(n2253), .A(n2250), .S(n6248), .Y(n2257) );
  MUX2X1 U5671 ( .B(n2256), .A(n2241), .S(n6233), .Y(n2259) );
  MUX2X1 U5672 ( .B(\Mem[62][1] ), .A(\Mem[63][1] ), .S(n6363), .Y(n2263) );
  MUX2X1 U5673 ( .B(\Mem[60][1] ), .A(\Mem[61][1] ), .S(n6363), .Y(n2262) );
  MUX2X1 U5674 ( .B(\Mem[58][1] ), .A(\Mem[59][1] ), .S(n6363), .Y(n2266) );
  MUX2X1 U5675 ( .B(\Mem[56][1] ), .A(\Mem[57][1] ), .S(n6363), .Y(n2265) );
  MUX2X1 U5676 ( .B(n2264), .A(n2261), .S(n6248), .Y(n2275) );
  MUX2X1 U5677 ( .B(\Mem[54][1] ), .A(\Mem[55][1] ), .S(n6364), .Y(n2269) );
  MUX2X1 U5678 ( .B(\Mem[52][1] ), .A(\Mem[53][1] ), .S(n6364), .Y(n2268) );
  MUX2X1 U5679 ( .B(\Mem[50][1] ), .A(\Mem[51][1] ), .S(n6364), .Y(n2272) );
  MUX2X1 U5680 ( .B(\Mem[48][1] ), .A(\Mem[49][1] ), .S(n6364), .Y(n2271) );
  MUX2X1 U5681 ( .B(n2270), .A(n2267), .S(n6249), .Y(n2274) );
  MUX2X1 U5682 ( .B(\Mem[46][1] ), .A(\Mem[47][1] ), .S(n6364), .Y(n2278) );
  MUX2X1 U5683 ( .B(\Mem[44][1] ), .A(\Mem[45][1] ), .S(n6364), .Y(n2277) );
  MUX2X1 U5684 ( .B(\Mem[42][1] ), .A(\Mem[43][1] ), .S(n6364), .Y(n2281) );
  MUX2X1 U5685 ( .B(\Mem[40][1] ), .A(\Mem[41][1] ), .S(n6364), .Y(n2280) );
  MUX2X1 U5686 ( .B(n2279), .A(n2276), .S(n6249), .Y(n4338) );
  MUX2X1 U5687 ( .B(\Mem[38][1] ), .A(\Mem[39][1] ), .S(n6364), .Y(n2284) );
  MUX2X1 U5688 ( .B(\Mem[36][1] ), .A(\Mem[37][1] ), .S(n6364), .Y(n2283) );
  MUX2X1 U5689 ( .B(\Mem[34][1] ), .A(\Mem[35][1] ), .S(n6364), .Y(n4335) );
  MUX2X1 U5690 ( .B(\Mem[32][1] ), .A(\Mem[33][1] ), .S(n6364), .Y(n4334) );
  MUX2X1 U5691 ( .B(n2285), .A(n2282), .S(n6249), .Y(n4337) );
  MUX2X1 U5692 ( .B(n4336), .A(n2273), .S(n6233), .Y(n4370) );
  MUX2X1 U5693 ( .B(\Mem[30][1] ), .A(\Mem[31][1] ), .S(n6364), .Y(n4341) );
  MUX2X1 U5694 ( .B(\Mem[28][1] ), .A(\Mem[29][1] ), .S(n6365), .Y(n4340) );
  MUX2X1 U5695 ( .B(\Mem[26][1] ), .A(\Mem[27][1] ), .S(n6365), .Y(n4344) );
  MUX2X1 U5696 ( .B(\Mem[24][1] ), .A(\Mem[25][1] ), .S(n6365), .Y(n4343) );
  MUX2X1 U5697 ( .B(n4342), .A(n4339), .S(n6249), .Y(n4353) );
  MUX2X1 U5698 ( .B(\Mem[22][1] ), .A(\Mem[23][1] ), .S(n6365), .Y(n4347) );
  MUX2X1 U5699 ( .B(\Mem[20][1] ), .A(\Mem[21][1] ), .S(n6365), .Y(n4346) );
  MUX2X1 U5700 ( .B(\Mem[18][1] ), .A(\Mem[19][1] ), .S(n6365), .Y(n4350) );
  MUX2X1 U5701 ( .B(\Mem[16][1] ), .A(\Mem[17][1] ), .S(n6365), .Y(n4349) );
  MUX2X1 U5702 ( .B(n4348), .A(n4345), .S(n6249), .Y(n4352) );
  MUX2X1 U5703 ( .B(\Mem[14][1] ), .A(\Mem[15][1] ), .S(n6365), .Y(n4356) );
  MUX2X1 U5704 ( .B(\Mem[12][1] ), .A(\Mem[13][1] ), .S(n6365), .Y(n4355) );
  MUX2X1 U5705 ( .B(\Mem[10][1] ), .A(\Mem[11][1] ), .S(n6365), .Y(n4359) );
  MUX2X1 U5706 ( .B(\Mem[8][1] ), .A(\Mem[9][1] ), .S(n6365), .Y(n4358) );
  MUX2X1 U5707 ( .B(n4357), .A(n4354), .S(n6249), .Y(n4368) );
  MUX2X1 U5708 ( .B(\Mem[6][1] ), .A(\Mem[7][1] ), .S(n6365), .Y(n4362) );
  MUX2X1 U5709 ( .B(\Mem[4][1] ), .A(\Mem[5][1] ), .S(n6365), .Y(n4361) );
  MUX2X1 U5710 ( .B(\Mem[2][1] ), .A(\Mem[3][1] ), .S(n6366), .Y(n4365) );
  MUX2X1 U5711 ( .B(\Mem[0][1] ), .A(\Mem[1][1] ), .S(n6366), .Y(n4364) );
  MUX2X1 U5712 ( .B(n4363), .A(n4360), .S(n6249), .Y(n4367) );
  MUX2X1 U5713 ( .B(n4366), .A(n4351), .S(n6233), .Y(n4369) );
  MUX2X1 U5714 ( .B(\Mem[62][2] ), .A(\Mem[63][2] ), .S(n6366), .Y(n4373) );
  MUX2X1 U5715 ( .B(\Mem[60][2] ), .A(\Mem[61][2] ), .S(n6366), .Y(n4372) );
  MUX2X1 U5716 ( .B(\Mem[58][2] ), .A(\Mem[59][2] ), .S(n6366), .Y(n4376) );
  MUX2X1 U5717 ( .B(\Mem[56][2] ), .A(\Mem[57][2] ), .S(n6366), .Y(n4375) );
  MUX2X1 U5718 ( .B(n4374), .A(n4371), .S(n6249), .Y(n4385) );
  MUX2X1 U5719 ( .B(\Mem[54][2] ), .A(\Mem[55][2] ), .S(n6366), .Y(n4379) );
  MUX2X1 U5720 ( .B(\Mem[52][2] ), .A(\Mem[53][2] ), .S(n6366), .Y(n4378) );
  MUX2X1 U5721 ( .B(\Mem[50][2] ), .A(\Mem[51][2] ), .S(n6366), .Y(n4382) );
  MUX2X1 U5722 ( .B(\Mem[48][2] ), .A(\Mem[49][2] ), .S(n6366), .Y(n4381) );
  MUX2X1 U5723 ( .B(n4380), .A(n4377), .S(n6249), .Y(n4384) );
  MUX2X1 U5724 ( .B(\Mem[46][2] ), .A(\Mem[47][2] ), .S(n6366), .Y(n4388) );
  MUX2X1 U5725 ( .B(\Mem[44][2] ), .A(\Mem[45][2] ), .S(n6366), .Y(n4387) );
  MUX2X1 U5726 ( .B(\Mem[42][2] ), .A(\Mem[43][2] ), .S(n6366), .Y(n4391) );
  MUX2X1 U5727 ( .B(\Mem[40][2] ), .A(\Mem[41][2] ), .S(n6367), .Y(n4390) );
  MUX2X1 U5728 ( .B(n4389), .A(n4386), .S(n6249), .Y(n4400) );
  MUX2X1 U5729 ( .B(\Mem[38][2] ), .A(\Mem[39][2] ), .S(n6367), .Y(n4394) );
  MUX2X1 U5730 ( .B(\Mem[36][2] ), .A(\Mem[37][2] ), .S(n6367), .Y(n4393) );
  MUX2X1 U5731 ( .B(\Mem[34][2] ), .A(\Mem[35][2] ), .S(n6367), .Y(n4397) );
  MUX2X1 U5732 ( .B(\Mem[32][2] ), .A(\Mem[33][2] ), .S(n6367), .Y(n4396) );
  MUX2X1 U5733 ( .B(n4395), .A(n4392), .S(n6249), .Y(n4399) );
  MUX2X1 U5734 ( .B(n4398), .A(n4383), .S(n6233), .Y(n4432) );
  MUX2X1 U5735 ( .B(\Mem[30][2] ), .A(\Mem[31][2] ), .S(n6367), .Y(n4403) );
  MUX2X1 U5736 ( .B(\Mem[28][2] ), .A(\Mem[29][2] ), .S(n6367), .Y(n4402) );
  MUX2X1 U5737 ( .B(\Mem[26][2] ), .A(\Mem[27][2] ), .S(n6367), .Y(n4406) );
  MUX2X1 U5738 ( .B(\Mem[24][2] ), .A(\Mem[25][2] ), .S(n6367), .Y(n4405) );
  MUX2X1 U5739 ( .B(n4404), .A(n4401), .S(n6249), .Y(n4415) );
  MUX2X1 U5740 ( .B(\Mem[22][2] ), .A(\Mem[23][2] ), .S(n6367), .Y(n4409) );
  MUX2X1 U5741 ( .B(\Mem[20][2] ), .A(\Mem[21][2] ), .S(n6367), .Y(n4408) );
  MUX2X1 U5742 ( .B(\Mem[18][2] ), .A(\Mem[19][2] ), .S(n6367), .Y(n4412) );
  MUX2X1 U5743 ( .B(\Mem[16][2] ), .A(\Mem[17][2] ), .S(n6367), .Y(n4411) );
  MUX2X1 U5744 ( .B(n4410), .A(n4407), .S(n6249), .Y(n4414) );
  MUX2X1 U5745 ( .B(\Mem[14][2] ), .A(\Mem[15][2] ), .S(n6368), .Y(n4418) );
  MUX2X1 U5746 ( .B(\Mem[12][2] ), .A(\Mem[13][2] ), .S(n6368), .Y(n4417) );
  MUX2X1 U5747 ( .B(\Mem[10][2] ), .A(\Mem[11][2] ), .S(n6368), .Y(n4421) );
  MUX2X1 U5748 ( .B(\Mem[8][2] ), .A(\Mem[9][2] ), .S(n6368), .Y(n4420) );
  MUX2X1 U5749 ( .B(n4419), .A(n4416), .S(n6250), .Y(n4430) );
  MUX2X1 U5750 ( .B(\Mem[6][2] ), .A(\Mem[7][2] ), .S(n6368), .Y(n4424) );
  MUX2X1 U5751 ( .B(\Mem[4][2] ), .A(\Mem[5][2] ), .S(n6368), .Y(n4423) );
  MUX2X1 U5752 ( .B(\Mem[2][2] ), .A(\Mem[3][2] ), .S(n6368), .Y(n4427) );
  MUX2X1 U5753 ( .B(\Mem[0][2] ), .A(\Mem[1][2] ), .S(n6368), .Y(n4426) );
  MUX2X1 U5754 ( .B(n4425), .A(n4422), .S(n6250), .Y(n4429) );
  MUX2X1 U5755 ( .B(n4428), .A(n4413), .S(n6233), .Y(n4431) );
  MUX2X1 U5756 ( .B(\Mem[62][3] ), .A(\Mem[63][3] ), .S(n6368), .Y(n4435) );
  MUX2X1 U5757 ( .B(\Mem[60][3] ), .A(\Mem[61][3] ), .S(n6368), .Y(n4434) );
  MUX2X1 U5758 ( .B(\Mem[58][3] ), .A(\Mem[59][3] ), .S(n6368), .Y(n4438) );
  MUX2X1 U5759 ( .B(\Mem[56][3] ), .A(\Mem[57][3] ), .S(n6368), .Y(n4437) );
  MUX2X1 U5760 ( .B(n4436), .A(n4433), .S(n6250), .Y(n4447) );
  MUX2X1 U5761 ( .B(\Mem[54][3] ), .A(\Mem[55][3] ), .S(n6368), .Y(n4441) );
  MUX2X1 U5762 ( .B(\Mem[52][3] ), .A(\Mem[53][3] ), .S(n6369), .Y(n4440) );
  MUX2X1 U5763 ( .B(\Mem[50][3] ), .A(\Mem[51][3] ), .S(n6369), .Y(n4444) );
  MUX2X1 U5764 ( .B(\Mem[48][3] ), .A(\Mem[49][3] ), .S(n6369), .Y(n4443) );
  MUX2X1 U5765 ( .B(n4442), .A(n4439), .S(n6250), .Y(n4446) );
  MUX2X1 U5766 ( .B(\Mem[46][3] ), .A(\Mem[47][3] ), .S(n6369), .Y(n4450) );
  MUX2X1 U5767 ( .B(\Mem[44][3] ), .A(\Mem[45][3] ), .S(n6369), .Y(n4449) );
  MUX2X1 U5768 ( .B(\Mem[42][3] ), .A(\Mem[43][3] ), .S(n6369), .Y(n4453) );
  MUX2X1 U5769 ( .B(\Mem[40][3] ), .A(\Mem[41][3] ), .S(n6369), .Y(n4452) );
  MUX2X1 U5770 ( .B(n4451), .A(n4448), .S(n6250), .Y(n4462) );
  MUX2X1 U5771 ( .B(\Mem[38][3] ), .A(\Mem[39][3] ), .S(n6369), .Y(n4456) );
  MUX2X1 U5772 ( .B(\Mem[36][3] ), .A(\Mem[37][3] ), .S(n6369), .Y(n4455) );
  MUX2X1 U5773 ( .B(\Mem[34][3] ), .A(\Mem[35][3] ), .S(n6369), .Y(n4459) );
  MUX2X1 U5774 ( .B(\Mem[32][3] ), .A(\Mem[33][3] ), .S(n6369), .Y(n4458) );
  MUX2X1 U5775 ( .B(n4457), .A(n4454), .S(n6250), .Y(n4461) );
  MUX2X1 U5776 ( .B(n4460), .A(n4445), .S(n6233), .Y(n4494) );
  MUX2X1 U5777 ( .B(\Mem[30][3] ), .A(\Mem[31][3] ), .S(n6369), .Y(n4465) );
  MUX2X1 U5778 ( .B(\Mem[28][3] ), .A(\Mem[29][3] ), .S(n6369), .Y(n4464) );
  MUX2X1 U5779 ( .B(\Mem[26][3] ), .A(\Mem[27][3] ), .S(n6370), .Y(n4468) );
  MUX2X1 U5780 ( .B(\Mem[24][3] ), .A(\Mem[25][3] ), .S(n6370), .Y(n4467) );
  MUX2X1 U5781 ( .B(n4466), .A(n4463), .S(n6250), .Y(n4477) );
  MUX2X1 U5782 ( .B(\Mem[22][3] ), .A(\Mem[23][3] ), .S(n6370), .Y(n4471) );
  MUX2X1 U5783 ( .B(\Mem[20][3] ), .A(\Mem[21][3] ), .S(n6370), .Y(n4470) );
  MUX2X1 U5784 ( .B(\Mem[18][3] ), .A(\Mem[19][3] ), .S(n6370), .Y(n4474) );
  MUX2X1 U5785 ( .B(\Mem[16][3] ), .A(\Mem[17][3] ), .S(n6370), .Y(n4473) );
  MUX2X1 U5786 ( .B(n4472), .A(n4469), .S(n6250), .Y(n4476) );
  MUX2X1 U5787 ( .B(\Mem[14][3] ), .A(\Mem[15][3] ), .S(n6370), .Y(n4480) );
  MUX2X1 U5788 ( .B(\Mem[12][3] ), .A(\Mem[13][3] ), .S(n6370), .Y(n4479) );
  MUX2X1 U5789 ( .B(\Mem[10][3] ), .A(\Mem[11][3] ), .S(n6370), .Y(n4483) );
  MUX2X1 U5790 ( .B(\Mem[8][3] ), .A(\Mem[9][3] ), .S(n6370), .Y(n4482) );
  MUX2X1 U5791 ( .B(n4481), .A(n4478), .S(n6250), .Y(n4492) );
  MUX2X1 U5792 ( .B(\Mem[6][3] ), .A(\Mem[7][3] ), .S(n6370), .Y(n4486) );
  MUX2X1 U5793 ( .B(\Mem[4][3] ), .A(\Mem[5][3] ), .S(n6370), .Y(n4485) );
  MUX2X1 U5794 ( .B(\Mem[2][3] ), .A(\Mem[3][3] ), .S(n6370), .Y(n4489) );
  MUX2X1 U5795 ( .B(\Mem[0][3] ), .A(\Mem[1][3] ), .S(n6371), .Y(n4488) );
  MUX2X1 U5796 ( .B(n4487), .A(n4484), .S(n6250), .Y(n4491) );
  MUX2X1 U5797 ( .B(n4490), .A(n4475), .S(n6233), .Y(n4493) );
  MUX2X1 U5798 ( .B(\Mem[62][4] ), .A(\Mem[63][4] ), .S(n6371), .Y(n4497) );
  MUX2X1 U5799 ( .B(\Mem[60][4] ), .A(\Mem[61][4] ), .S(n6371), .Y(n4496) );
  MUX2X1 U5800 ( .B(\Mem[58][4] ), .A(\Mem[59][4] ), .S(n6371), .Y(n4500) );
  MUX2X1 U5801 ( .B(\Mem[56][4] ), .A(\Mem[57][4] ), .S(n6371), .Y(n4499) );
  MUX2X1 U5802 ( .B(n4498), .A(n4495), .S(n6250), .Y(n4509) );
  MUX2X1 U5803 ( .B(\Mem[54][4] ), .A(\Mem[55][4] ), .S(n6371), .Y(n4503) );
  MUX2X1 U5804 ( .B(\Mem[52][4] ), .A(\Mem[53][4] ), .S(n6371), .Y(n4502) );
  MUX2X1 U5805 ( .B(\Mem[50][4] ), .A(\Mem[51][4] ), .S(n6371), .Y(n4506) );
  MUX2X1 U5806 ( .B(\Mem[48][4] ), .A(\Mem[49][4] ), .S(n6371), .Y(n4505) );
  MUX2X1 U5807 ( .B(n4504), .A(n4501), .S(n6250), .Y(n4508) );
  MUX2X1 U5808 ( .B(\Mem[46][4] ), .A(\Mem[47][4] ), .S(n6371), .Y(n4512) );
  MUX2X1 U5809 ( .B(\Mem[44][4] ), .A(\Mem[45][4] ), .S(n6371), .Y(n4511) );
  MUX2X1 U5810 ( .B(\Mem[42][4] ), .A(\Mem[43][4] ), .S(n6371), .Y(n4515) );
  MUX2X1 U5811 ( .B(\Mem[40][4] ), .A(\Mem[41][4] ), .S(n6371), .Y(n4514) );
  MUX2X1 U5812 ( .B(n4513), .A(n4510), .S(n6250), .Y(n4524) );
  MUX2X1 U5813 ( .B(\Mem[38][4] ), .A(\Mem[39][4] ), .S(n6372), .Y(n4518) );
  MUX2X1 U5814 ( .B(\Mem[36][4] ), .A(\Mem[37][4] ), .S(n6372), .Y(n4517) );
  MUX2X1 U5815 ( .B(\Mem[34][4] ), .A(\Mem[35][4] ), .S(n6372), .Y(n4521) );
  MUX2X1 U5816 ( .B(\Mem[32][4] ), .A(\Mem[33][4] ), .S(n6372), .Y(n4520) );
  MUX2X1 U5817 ( .B(n4519), .A(n4516), .S(n6251), .Y(n4523) );
  MUX2X1 U5818 ( .B(n4522), .A(n4507), .S(n6233), .Y(n4556) );
  MUX2X1 U5819 ( .B(\Mem[30][4] ), .A(\Mem[31][4] ), .S(n6372), .Y(n4527) );
  MUX2X1 U5820 ( .B(\Mem[28][4] ), .A(\Mem[29][4] ), .S(n6372), .Y(n4526) );
  MUX2X1 U5821 ( .B(\Mem[26][4] ), .A(\Mem[27][4] ), .S(n6372), .Y(n4530) );
  MUX2X1 U5822 ( .B(\Mem[24][4] ), .A(\Mem[25][4] ), .S(n6372), .Y(n4529) );
  MUX2X1 U5823 ( .B(n4528), .A(n4525), .S(n6251), .Y(n4539) );
  MUX2X1 U5824 ( .B(\Mem[22][4] ), .A(\Mem[23][4] ), .S(n6372), .Y(n4533) );
  MUX2X1 U5825 ( .B(\Mem[20][4] ), .A(\Mem[21][4] ), .S(n6372), .Y(n4532) );
  MUX2X1 U5826 ( .B(\Mem[18][4] ), .A(\Mem[19][4] ), .S(n6372), .Y(n4536) );
  MUX2X1 U5827 ( .B(\Mem[16][4] ), .A(\Mem[17][4] ), .S(n6372), .Y(n4535) );
  MUX2X1 U5828 ( .B(n4534), .A(n4531), .S(n6251), .Y(n4538) );
  MUX2X1 U5829 ( .B(\Mem[14][4] ), .A(\Mem[15][4] ), .S(n6372), .Y(n4542) );
  MUX2X1 U5830 ( .B(\Mem[12][4] ), .A(\Mem[13][4] ), .S(n6373), .Y(n4541) );
  MUX2X1 U5831 ( .B(\Mem[10][4] ), .A(\Mem[11][4] ), .S(n6373), .Y(n4545) );
  MUX2X1 U5832 ( .B(\Mem[8][4] ), .A(\Mem[9][4] ), .S(n6373), .Y(n4544) );
  MUX2X1 U5833 ( .B(n4543), .A(n4540), .S(n6251), .Y(n4554) );
  MUX2X1 U5834 ( .B(\Mem[6][4] ), .A(\Mem[7][4] ), .S(n6373), .Y(n4548) );
  MUX2X1 U5835 ( .B(\Mem[4][4] ), .A(\Mem[5][4] ), .S(n6373), .Y(n4547) );
  MUX2X1 U5836 ( .B(\Mem[2][4] ), .A(\Mem[3][4] ), .S(n6373), .Y(n4551) );
  MUX2X1 U5837 ( .B(\Mem[0][4] ), .A(\Mem[1][4] ), .S(n6373), .Y(n4550) );
  MUX2X1 U5838 ( .B(n4549), .A(n4546), .S(n6251), .Y(n4553) );
  MUX2X1 U5839 ( .B(n4552), .A(n4537), .S(n6233), .Y(n4555) );
  MUX2X1 U5840 ( .B(\Mem[62][5] ), .A(\Mem[63][5] ), .S(n6373), .Y(n4559) );
  MUX2X1 U5841 ( .B(\Mem[60][5] ), .A(\Mem[61][5] ), .S(n6373), .Y(n4558) );
  MUX2X1 U5842 ( .B(\Mem[58][5] ), .A(\Mem[59][5] ), .S(n6373), .Y(n4562) );
  MUX2X1 U5843 ( .B(\Mem[56][5] ), .A(\Mem[57][5] ), .S(n6373), .Y(n4561) );
  MUX2X1 U5844 ( .B(n4560), .A(n4557), .S(n6251), .Y(n4571) );
  MUX2X1 U5845 ( .B(\Mem[54][5] ), .A(\Mem[55][5] ), .S(n6373), .Y(n4565) );
  MUX2X1 U5846 ( .B(\Mem[52][5] ), .A(\Mem[53][5] ), .S(n6373), .Y(n4564) );
  MUX2X1 U5847 ( .B(\Mem[50][5] ), .A(\Mem[51][5] ), .S(n6374), .Y(n4568) );
  MUX2X1 U5848 ( .B(\Mem[48][5] ), .A(\Mem[49][5] ), .S(n6374), .Y(n4567) );
  MUX2X1 U5849 ( .B(n4566), .A(n4563), .S(n6251), .Y(n4570) );
  MUX2X1 U5850 ( .B(\Mem[46][5] ), .A(\Mem[47][5] ), .S(n6374), .Y(n4574) );
  MUX2X1 U5851 ( .B(\Mem[44][5] ), .A(\Mem[45][5] ), .S(n6374), .Y(n4573) );
  MUX2X1 U5852 ( .B(\Mem[42][5] ), .A(\Mem[43][5] ), .S(n6374), .Y(n4577) );
  MUX2X1 U5853 ( .B(\Mem[40][5] ), .A(\Mem[41][5] ), .S(n6374), .Y(n4576) );
  MUX2X1 U5854 ( .B(n4575), .A(n4572), .S(n6251), .Y(n4586) );
  MUX2X1 U5855 ( .B(\Mem[38][5] ), .A(\Mem[39][5] ), .S(n6374), .Y(n4580) );
  MUX2X1 U5856 ( .B(\Mem[36][5] ), .A(\Mem[37][5] ), .S(n6374), .Y(n4579) );
  MUX2X1 U5857 ( .B(\Mem[34][5] ), .A(\Mem[35][5] ), .S(n6374), .Y(n4583) );
  MUX2X1 U5858 ( .B(\Mem[32][5] ), .A(\Mem[33][5] ), .S(n6374), .Y(n4582) );
  MUX2X1 U5859 ( .B(n4581), .A(n4578), .S(n6251), .Y(n4585) );
  MUX2X1 U5860 ( .B(n4584), .A(n4569), .S(n6233), .Y(n4618) );
  MUX2X1 U5861 ( .B(\Mem[30][5] ), .A(\Mem[31][5] ), .S(n6374), .Y(n4589) );
  MUX2X1 U5862 ( .B(\Mem[28][5] ), .A(\Mem[29][5] ), .S(n6374), .Y(n4588) );
  MUX2X1 U5863 ( .B(\Mem[26][5] ), .A(\Mem[27][5] ), .S(n6374), .Y(n4592) );
  MUX2X1 U5864 ( .B(\Mem[24][5] ), .A(\Mem[25][5] ), .S(n6375), .Y(n4591) );
  MUX2X1 U5865 ( .B(n4590), .A(n4587), .S(n6251), .Y(n4601) );
  MUX2X1 U5866 ( .B(\Mem[22][5] ), .A(\Mem[23][5] ), .S(n6375), .Y(n4595) );
  MUX2X1 U5867 ( .B(\Mem[20][5] ), .A(\Mem[21][5] ), .S(n6375), .Y(n4594) );
  MUX2X1 U5868 ( .B(\Mem[18][5] ), .A(\Mem[19][5] ), .S(n6375), .Y(n4598) );
  MUX2X1 U5869 ( .B(\Mem[16][5] ), .A(\Mem[17][5] ), .S(n6375), .Y(n4597) );
  MUX2X1 U5870 ( .B(n4596), .A(n4593), .S(n6251), .Y(n4600) );
  MUX2X1 U5871 ( .B(\Mem[14][5] ), .A(\Mem[15][5] ), .S(n6375), .Y(n4604) );
  MUX2X1 U5872 ( .B(\Mem[12][5] ), .A(\Mem[13][5] ), .S(n6375), .Y(n4603) );
  MUX2X1 U5873 ( .B(\Mem[10][5] ), .A(\Mem[11][5] ), .S(n6375), .Y(n4607) );
  MUX2X1 U5874 ( .B(\Mem[8][5] ), .A(\Mem[9][5] ), .S(n6375), .Y(n4606) );
  MUX2X1 U5875 ( .B(n4605), .A(n4602), .S(n6251), .Y(n4616) );
  MUX2X1 U5876 ( .B(\Mem[6][5] ), .A(\Mem[7][5] ), .S(n6375), .Y(n4610) );
  MUX2X1 U5877 ( .B(\Mem[4][5] ), .A(\Mem[5][5] ), .S(n6375), .Y(n4609) );
  MUX2X1 U5878 ( .B(\Mem[2][5] ), .A(\Mem[3][5] ), .S(n6375), .Y(n4613) );
  MUX2X1 U5879 ( .B(\Mem[0][5] ), .A(\Mem[1][5] ), .S(n6375), .Y(n4612) );
  MUX2X1 U5880 ( .B(n4611), .A(n4608), .S(n6251), .Y(n4615) );
  MUX2X1 U5881 ( .B(n4614), .A(n4599), .S(n6233), .Y(n4617) );
  MUX2X1 U5882 ( .B(\Mem[62][6] ), .A(\Mem[63][6] ), .S(n6376), .Y(n4621) );
  MUX2X1 U5883 ( .B(\Mem[60][6] ), .A(\Mem[61][6] ), .S(n6376), .Y(n4620) );
  MUX2X1 U5884 ( .B(\Mem[58][6] ), .A(\Mem[59][6] ), .S(n6376), .Y(n4624) );
  MUX2X1 U5885 ( .B(\Mem[56][6] ), .A(\Mem[57][6] ), .S(n6376), .Y(n4623) );
  MUX2X1 U5886 ( .B(n4622), .A(n4619), .S(n6252), .Y(n4633) );
  MUX2X1 U5887 ( .B(\Mem[54][6] ), .A(\Mem[55][6] ), .S(n6376), .Y(n4627) );
  MUX2X1 U5888 ( .B(\Mem[52][6] ), .A(\Mem[53][6] ), .S(n6376), .Y(n4626) );
  MUX2X1 U5889 ( .B(\Mem[50][6] ), .A(\Mem[51][6] ), .S(n6376), .Y(n4630) );
  MUX2X1 U5890 ( .B(\Mem[48][6] ), .A(\Mem[49][6] ), .S(n6376), .Y(n4629) );
  MUX2X1 U5891 ( .B(n4628), .A(n4625), .S(n6252), .Y(n4632) );
  MUX2X1 U5892 ( .B(\Mem[46][6] ), .A(\Mem[47][6] ), .S(n6376), .Y(n4636) );
  MUX2X1 U5893 ( .B(\Mem[44][6] ), .A(\Mem[45][6] ), .S(n6376), .Y(n4635) );
  MUX2X1 U5894 ( .B(\Mem[42][6] ), .A(\Mem[43][6] ), .S(n6376), .Y(n4639) );
  MUX2X1 U5895 ( .B(\Mem[40][6] ), .A(\Mem[41][6] ), .S(n6376), .Y(n4638) );
  MUX2X1 U5896 ( .B(n4637), .A(n4634), .S(n6252), .Y(n4648) );
  MUX2X1 U5897 ( .B(\Mem[38][6] ), .A(\Mem[39][6] ), .S(n6376), .Y(n4642) );
  MUX2X1 U5898 ( .B(\Mem[36][6] ), .A(\Mem[37][6] ), .S(n6377), .Y(n4641) );
  MUX2X1 U5899 ( .B(\Mem[34][6] ), .A(\Mem[35][6] ), .S(n6377), .Y(n4645) );
  MUX2X1 U5900 ( .B(\Mem[32][6] ), .A(\Mem[33][6] ), .S(n6377), .Y(n4644) );
  MUX2X1 U5901 ( .B(n4643), .A(n4640), .S(n6252), .Y(n4647) );
  MUX2X1 U5902 ( .B(n4646), .A(n4631), .S(n6234), .Y(n4680) );
  MUX2X1 U5903 ( .B(\Mem[30][6] ), .A(\Mem[31][6] ), .S(n6377), .Y(n4651) );
  MUX2X1 U5904 ( .B(\Mem[28][6] ), .A(\Mem[29][6] ), .S(n6377), .Y(n4650) );
  MUX2X1 U5905 ( .B(\Mem[26][6] ), .A(\Mem[27][6] ), .S(n6377), .Y(n4654) );
  MUX2X1 U5906 ( .B(\Mem[24][6] ), .A(\Mem[25][6] ), .S(n6377), .Y(n4653) );
  MUX2X1 U5907 ( .B(n4652), .A(n4649), .S(n6252), .Y(n4663) );
  MUX2X1 U5908 ( .B(\Mem[22][6] ), .A(\Mem[23][6] ), .S(n6377), .Y(n4657) );
  MUX2X1 U5909 ( .B(\Mem[20][6] ), .A(\Mem[21][6] ), .S(n6377), .Y(n4656) );
  MUX2X1 U5910 ( .B(\Mem[18][6] ), .A(\Mem[19][6] ), .S(n6377), .Y(n4660) );
  MUX2X1 U5911 ( .B(\Mem[16][6] ), .A(\Mem[17][6] ), .S(n6377), .Y(n4659) );
  MUX2X1 U5912 ( .B(n4658), .A(n4655), .S(n6252), .Y(n4662) );
  MUX2X1 U5913 ( .B(\Mem[14][6] ), .A(\Mem[15][6] ), .S(n6377), .Y(n4666) );
  MUX2X1 U5914 ( .B(\Mem[12][6] ), .A(\Mem[13][6] ), .S(n6377), .Y(n4665) );
  MUX2X1 U5915 ( .B(\Mem[10][6] ), .A(\Mem[11][6] ), .S(n6378), .Y(n4669) );
  MUX2X1 U5916 ( .B(\Mem[8][6] ), .A(\Mem[9][6] ), .S(n6378), .Y(n4668) );
  MUX2X1 U5917 ( .B(n4667), .A(n4664), .S(n6252), .Y(n4678) );
  MUX2X1 U5918 ( .B(\Mem[6][6] ), .A(\Mem[7][6] ), .S(n6378), .Y(n4672) );
  MUX2X1 U5919 ( .B(\Mem[4][6] ), .A(\Mem[5][6] ), .S(n6378), .Y(n4671) );
  MUX2X1 U5920 ( .B(\Mem[2][6] ), .A(\Mem[3][6] ), .S(n6378), .Y(n4675) );
  MUX2X1 U5921 ( .B(\Mem[0][6] ), .A(\Mem[1][6] ), .S(n6378), .Y(n4674) );
  MUX2X1 U5922 ( .B(n4673), .A(n4670), .S(n6252), .Y(n4677) );
  MUX2X1 U5923 ( .B(n4676), .A(n4661), .S(n6234), .Y(n4679) );
  MUX2X1 U5924 ( .B(\Mem[62][7] ), .A(\Mem[63][7] ), .S(n6378), .Y(n4683) );
  MUX2X1 U5925 ( .B(\Mem[60][7] ), .A(\Mem[61][7] ), .S(n6378), .Y(n4682) );
  MUX2X1 U5926 ( .B(\Mem[58][7] ), .A(\Mem[59][7] ), .S(n6378), .Y(n4686) );
  MUX2X1 U5927 ( .B(\Mem[56][7] ), .A(\Mem[57][7] ), .S(n6378), .Y(n4685) );
  MUX2X1 U5928 ( .B(n4684), .A(n4681), .S(n6252), .Y(n4695) );
  MUX2X1 U5929 ( .B(\Mem[54][7] ), .A(\Mem[55][7] ), .S(n6378), .Y(n4689) );
  MUX2X1 U5930 ( .B(\Mem[52][7] ), .A(\Mem[53][7] ), .S(n6378), .Y(n4688) );
  MUX2X1 U5931 ( .B(\Mem[50][7] ), .A(\Mem[51][7] ), .S(n6378), .Y(n4692) );
  MUX2X1 U5932 ( .B(\Mem[48][7] ), .A(\Mem[49][7] ), .S(n6379), .Y(n4691) );
  MUX2X1 U5933 ( .B(n4690), .A(n4687), .S(n6252), .Y(n4694) );
  MUX2X1 U5934 ( .B(\Mem[46][7] ), .A(\Mem[47][7] ), .S(n6379), .Y(n4698) );
  MUX2X1 U5935 ( .B(\Mem[44][7] ), .A(\Mem[45][7] ), .S(n6379), .Y(n4697) );
  MUX2X1 U5936 ( .B(\Mem[42][7] ), .A(\Mem[43][7] ), .S(n6379), .Y(n4701) );
  MUX2X1 U5937 ( .B(\Mem[40][7] ), .A(\Mem[41][7] ), .S(n6379), .Y(n4700) );
  MUX2X1 U5938 ( .B(n4699), .A(n4696), .S(n6252), .Y(n4710) );
  MUX2X1 U5939 ( .B(\Mem[38][7] ), .A(\Mem[39][7] ), .S(n6379), .Y(n4704) );
  MUX2X1 U5940 ( .B(\Mem[36][7] ), .A(\Mem[37][7] ), .S(n6379), .Y(n4703) );
  MUX2X1 U5941 ( .B(\Mem[34][7] ), .A(\Mem[35][7] ), .S(n6379), .Y(n4707) );
  MUX2X1 U5942 ( .B(\Mem[32][7] ), .A(\Mem[33][7] ), .S(n6379), .Y(n4706) );
  MUX2X1 U5943 ( .B(n4705), .A(n4702), .S(n6252), .Y(n4709) );
  MUX2X1 U5944 ( .B(n4708), .A(n4693), .S(n6234), .Y(n4742) );
  MUX2X1 U5945 ( .B(\Mem[30][7] ), .A(\Mem[31][7] ), .S(n6379), .Y(n4713) );
  MUX2X1 U5946 ( .B(\Mem[28][7] ), .A(\Mem[29][7] ), .S(n6379), .Y(n4712) );
  MUX2X1 U5947 ( .B(\Mem[26][7] ), .A(\Mem[27][7] ), .S(n6379), .Y(n4716) );
  MUX2X1 U5948 ( .B(\Mem[24][7] ), .A(\Mem[25][7] ), .S(n6379), .Y(n4715) );
  MUX2X1 U5949 ( .B(n4714), .A(n4711), .S(n6252), .Y(n4725) );
  MUX2X1 U5950 ( .B(\Mem[22][7] ), .A(\Mem[23][7] ), .S(n6380), .Y(n4719) );
  MUX2X1 U5951 ( .B(\Mem[20][7] ), .A(\Mem[21][7] ), .S(n6380), .Y(n4718) );
  MUX2X1 U5952 ( .B(\Mem[18][7] ), .A(\Mem[19][7] ), .S(n6380), .Y(n4722) );
  MUX2X1 U5953 ( .B(\Mem[16][7] ), .A(\Mem[17][7] ), .S(n6380), .Y(n4721) );
  MUX2X1 U5954 ( .B(n4720), .A(n4717), .S(n6253), .Y(n4724) );
  MUX2X1 U5955 ( .B(\Mem[14][7] ), .A(\Mem[15][7] ), .S(n6380), .Y(n4728) );
  MUX2X1 U5956 ( .B(\Mem[12][7] ), .A(\Mem[13][7] ), .S(n6380), .Y(n4727) );
  MUX2X1 U5957 ( .B(\Mem[10][7] ), .A(\Mem[11][7] ), .S(n6380), .Y(n4731) );
  MUX2X1 U5958 ( .B(\Mem[8][7] ), .A(\Mem[9][7] ), .S(n6380), .Y(n4730) );
  MUX2X1 U5959 ( .B(n4729), .A(n4726), .S(n6253), .Y(n4740) );
  MUX2X1 U5960 ( .B(\Mem[6][7] ), .A(\Mem[7][7] ), .S(n6380), .Y(n4734) );
  MUX2X1 U5961 ( .B(\Mem[4][7] ), .A(\Mem[5][7] ), .S(n6380), .Y(n4733) );
  MUX2X1 U5962 ( .B(\Mem[2][7] ), .A(\Mem[3][7] ), .S(n6380), .Y(n4737) );
  MUX2X1 U5963 ( .B(\Mem[0][7] ), .A(\Mem[1][7] ), .S(n6380), .Y(n4736) );
  MUX2X1 U5964 ( .B(n4735), .A(n4732), .S(n6253), .Y(n4739) );
  MUX2X1 U5965 ( .B(n4738), .A(n4723), .S(n6234), .Y(n4741) );
  MUX2X1 U5966 ( .B(\Mem[62][8] ), .A(\Mem[63][8] ), .S(n6380), .Y(n4745) );
  MUX2X1 U5967 ( .B(\Mem[60][8] ), .A(\Mem[61][8] ), .S(n6381), .Y(n4744) );
  MUX2X1 U5968 ( .B(\Mem[58][8] ), .A(\Mem[59][8] ), .S(n6381), .Y(n4748) );
  MUX2X1 U5969 ( .B(\Mem[56][8] ), .A(\Mem[57][8] ), .S(n6381), .Y(n4747) );
  MUX2X1 U5970 ( .B(n4746), .A(n4743), .S(n6253), .Y(n4757) );
  MUX2X1 U5971 ( .B(\Mem[54][8] ), .A(\Mem[55][8] ), .S(n6381), .Y(n4751) );
  MUX2X1 U5972 ( .B(\Mem[52][8] ), .A(\Mem[53][8] ), .S(n6381), .Y(n4750) );
  MUX2X1 U5973 ( .B(\Mem[50][8] ), .A(\Mem[51][8] ), .S(n6381), .Y(n4754) );
  MUX2X1 U5974 ( .B(\Mem[48][8] ), .A(\Mem[49][8] ), .S(n6381), .Y(n4753) );
  MUX2X1 U5975 ( .B(n4752), .A(n4749), .S(n6253), .Y(n4756) );
  MUX2X1 U5976 ( .B(\Mem[46][8] ), .A(\Mem[47][8] ), .S(n6381), .Y(n4760) );
  MUX2X1 U5977 ( .B(\Mem[44][8] ), .A(\Mem[45][8] ), .S(n6381), .Y(n4759) );
  MUX2X1 U5978 ( .B(\Mem[42][8] ), .A(\Mem[43][8] ), .S(n6381), .Y(n4763) );
  MUX2X1 U5979 ( .B(\Mem[40][8] ), .A(\Mem[41][8] ), .S(n6381), .Y(n4762) );
  MUX2X1 U5980 ( .B(n4761), .A(n4758), .S(n6253), .Y(n4772) );
  MUX2X1 U5981 ( .B(\Mem[38][8] ), .A(\Mem[39][8] ), .S(n6381), .Y(n4766) );
  MUX2X1 U5982 ( .B(\Mem[36][8] ), .A(\Mem[37][8] ), .S(n6381), .Y(n4765) );
  MUX2X1 U5983 ( .B(\Mem[34][8] ), .A(\Mem[35][8] ), .S(n6382), .Y(n4769) );
  MUX2X1 U5984 ( .B(\Mem[32][8] ), .A(\Mem[33][8] ), .S(n6382), .Y(n4768) );
  MUX2X1 U5985 ( .B(n4767), .A(n4764), .S(n6253), .Y(n4771) );
  MUX2X1 U5986 ( .B(n4770), .A(n4755), .S(n6234), .Y(n4804) );
  MUX2X1 U5987 ( .B(\Mem[30][8] ), .A(\Mem[31][8] ), .S(n6382), .Y(n4775) );
  MUX2X1 U5988 ( .B(\Mem[28][8] ), .A(\Mem[29][8] ), .S(n6382), .Y(n4774) );
  MUX2X1 U5989 ( .B(\Mem[26][8] ), .A(\Mem[27][8] ), .S(n6382), .Y(n4778) );
  MUX2X1 U5990 ( .B(\Mem[24][8] ), .A(\Mem[25][8] ), .S(n6382), .Y(n4777) );
  MUX2X1 U5991 ( .B(n4776), .A(n4773), .S(n6253), .Y(n4787) );
  MUX2X1 U5992 ( .B(\Mem[22][8] ), .A(\Mem[23][8] ), .S(n6382), .Y(n4781) );
  MUX2X1 U5993 ( .B(\Mem[20][8] ), .A(\Mem[21][8] ), .S(n6382), .Y(n4780) );
  MUX2X1 U5994 ( .B(\Mem[18][8] ), .A(\Mem[19][8] ), .S(n6382), .Y(n4784) );
  MUX2X1 U5995 ( .B(\Mem[16][8] ), .A(\Mem[17][8] ), .S(n6382), .Y(n4783) );
  MUX2X1 U5996 ( .B(n4782), .A(n4779), .S(n6253), .Y(n4786) );
  MUX2X1 U5997 ( .B(\Mem[14][8] ), .A(\Mem[15][8] ), .S(n6382), .Y(n4790) );
  MUX2X1 U5998 ( .B(\Mem[12][8] ), .A(\Mem[13][8] ), .S(n6382), .Y(n4789) );
  MUX2X1 U5999 ( .B(\Mem[10][8] ), .A(\Mem[11][8] ), .S(n6382), .Y(n4793) );
  MUX2X1 U6000 ( .B(\Mem[8][8] ), .A(\Mem[9][8] ), .S(n6383), .Y(n4792) );
  MUX2X1 U6001 ( .B(n4791), .A(n4788), .S(n6253), .Y(n4802) );
  MUX2X1 U6002 ( .B(\Mem[6][8] ), .A(\Mem[7][8] ), .S(n6383), .Y(n4796) );
  MUX2X1 U6003 ( .B(\Mem[4][8] ), .A(\Mem[5][8] ), .S(n6383), .Y(n4795) );
  MUX2X1 U6004 ( .B(\Mem[2][8] ), .A(\Mem[3][8] ), .S(n6383), .Y(n4799) );
  MUX2X1 U6005 ( .B(\Mem[0][8] ), .A(\Mem[1][8] ), .S(n6383), .Y(n4798) );
  MUX2X1 U6006 ( .B(n4797), .A(n4794), .S(n6253), .Y(n4801) );
  MUX2X1 U6007 ( .B(n4800), .A(n4785), .S(n6234), .Y(n4803) );
  MUX2X1 U6008 ( .B(\Mem[62][9] ), .A(\Mem[63][9] ), .S(n6383), .Y(n4807) );
  MUX2X1 U6009 ( .B(\Mem[60][9] ), .A(\Mem[61][9] ), .S(n6383), .Y(n4806) );
  MUX2X1 U6010 ( .B(\Mem[58][9] ), .A(\Mem[59][9] ), .S(n6383), .Y(n4810) );
  MUX2X1 U6011 ( .B(\Mem[56][9] ), .A(\Mem[57][9] ), .S(n6383), .Y(n4809) );
  MUX2X1 U6012 ( .B(n4808), .A(n4805), .S(n6253), .Y(n4819) );
  MUX2X1 U6013 ( .B(\Mem[54][9] ), .A(\Mem[55][9] ), .S(n6383), .Y(n4813) );
  MUX2X1 U6014 ( .B(\Mem[52][9] ), .A(\Mem[53][9] ), .S(n6383), .Y(n4812) );
  MUX2X1 U6015 ( .B(\Mem[50][9] ), .A(\Mem[51][9] ), .S(n6383), .Y(n4816) );
  MUX2X1 U6016 ( .B(\Mem[48][9] ), .A(\Mem[49][9] ), .S(n6383), .Y(n4815) );
  MUX2X1 U6017 ( .B(n4814), .A(n4811), .S(n6253), .Y(n4818) );
  MUX2X1 U6018 ( .B(\Mem[46][9] ), .A(\Mem[47][9] ), .S(n6384), .Y(n4822) );
  MUX2X1 U6019 ( .B(\Mem[44][9] ), .A(\Mem[45][9] ), .S(n6384), .Y(n4821) );
  MUX2X1 U6020 ( .B(\Mem[42][9] ), .A(\Mem[43][9] ), .S(n6384), .Y(n4825) );
  MUX2X1 U6021 ( .B(\Mem[40][9] ), .A(\Mem[41][9] ), .S(n6384), .Y(n4824) );
  MUX2X1 U6022 ( .B(n4823), .A(n4820), .S(n6254), .Y(n4834) );
  MUX2X1 U6023 ( .B(\Mem[38][9] ), .A(\Mem[39][9] ), .S(n6384), .Y(n4828) );
  MUX2X1 U6024 ( .B(\Mem[36][9] ), .A(\Mem[37][9] ), .S(n6384), .Y(n4827) );
  MUX2X1 U6025 ( .B(\Mem[34][9] ), .A(\Mem[35][9] ), .S(n6384), .Y(n4831) );
  MUX2X1 U6026 ( .B(\Mem[32][9] ), .A(\Mem[33][9] ), .S(n6384), .Y(n4830) );
  MUX2X1 U6027 ( .B(n4829), .A(n4826), .S(n6254), .Y(n4833) );
  MUX2X1 U6028 ( .B(n4832), .A(n4817), .S(n6234), .Y(n4866) );
  MUX2X1 U6029 ( .B(\Mem[30][9] ), .A(\Mem[31][9] ), .S(n6384), .Y(n4837) );
  MUX2X1 U6030 ( .B(\Mem[28][9] ), .A(\Mem[29][9] ), .S(n6384), .Y(n4836) );
  MUX2X1 U6031 ( .B(\Mem[26][9] ), .A(\Mem[27][9] ), .S(n6384), .Y(n4840) );
  MUX2X1 U6032 ( .B(\Mem[24][9] ), .A(\Mem[25][9] ), .S(n6384), .Y(n4839) );
  MUX2X1 U6033 ( .B(n4838), .A(n4835), .S(n6254), .Y(n4849) );
  MUX2X1 U6034 ( .B(\Mem[22][9] ), .A(\Mem[23][9] ), .S(n6384), .Y(n4843) );
  MUX2X1 U6035 ( .B(\Mem[20][9] ), .A(\Mem[21][9] ), .S(n6385), .Y(n4842) );
  MUX2X1 U6036 ( .B(\Mem[18][9] ), .A(\Mem[19][9] ), .S(n6385), .Y(n4846) );
  MUX2X1 U6037 ( .B(\Mem[16][9] ), .A(\Mem[17][9] ), .S(n6385), .Y(n4845) );
  MUX2X1 U6038 ( .B(n4844), .A(n4841), .S(n6254), .Y(n4848) );
  MUX2X1 U6039 ( .B(\Mem[14][9] ), .A(\Mem[15][9] ), .S(n6385), .Y(n4852) );
  MUX2X1 U6040 ( .B(\Mem[12][9] ), .A(\Mem[13][9] ), .S(n6385), .Y(n4851) );
  MUX2X1 U6041 ( .B(\Mem[10][9] ), .A(\Mem[11][9] ), .S(n6385), .Y(n4855) );
  MUX2X1 U6042 ( .B(\Mem[8][9] ), .A(\Mem[9][9] ), .S(n6385), .Y(n4854) );
  MUX2X1 U6043 ( .B(n4853), .A(n4850), .S(n6254), .Y(n4864) );
  MUX2X1 U6044 ( .B(\Mem[6][9] ), .A(\Mem[7][9] ), .S(n6385), .Y(n4858) );
  MUX2X1 U6045 ( .B(\Mem[4][9] ), .A(\Mem[5][9] ), .S(n6385), .Y(n4857) );
  MUX2X1 U6046 ( .B(\Mem[2][9] ), .A(\Mem[3][9] ), .S(n6385), .Y(n4861) );
  MUX2X1 U6047 ( .B(\Mem[0][9] ), .A(\Mem[1][9] ), .S(n6385), .Y(n4860) );
  MUX2X1 U6048 ( .B(n4859), .A(n4856), .S(n6254), .Y(n4863) );
  MUX2X1 U6049 ( .B(n4862), .A(n4847), .S(n6234), .Y(n4865) );
  MUX2X1 U6050 ( .B(\Mem[62][10] ), .A(\Mem[63][10] ), .S(n6385), .Y(n4869) );
  MUX2X1 U6051 ( .B(\Mem[60][10] ), .A(\Mem[61][10] ), .S(n6385), .Y(n4868) );
  MUX2X1 U6052 ( .B(\Mem[58][10] ), .A(\Mem[59][10] ), .S(n6386), .Y(n4872) );
  MUX2X1 U6053 ( .B(\Mem[56][10] ), .A(\Mem[57][10] ), .S(n6386), .Y(n4871) );
  MUX2X1 U6054 ( .B(n4870), .A(n4867), .S(n6254), .Y(n4881) );
  MUX2X1 U6055 ( .B(\Mem[54][10] ), .A(\Mem[55][10] ), .S(n6386), .Y(n4875) );
  MUX2X1 U6056 ( .B(\Mem[52][10] ), .A(\Mem[53][10] ), .S(n6386), .Y(n4874) );
  MUX2X1 U6057 ( .B(\Mem[50][10] ), .A(\Mem[51][10] ), .S(n6386), .Y(n4878) );
  MUX2X1 U6058 ( .B(\Mem[48][10] ), .A(\Mem[49][10] ), .S(n6386), .Y(n4877) );
  MUX2X1 U6059 ( .B(n4876), .A(n4873), .S(n6254), .Y(n4880) );
  MUX2X1 U6060 ( .B(\Mem[46][10] ), .A(\Mem[47][10] ), .S(n6386), .Y(n4884) );
  MUX2X1 U6061 ( .B(\Mem[44][10] ), .A(\Mem[45][10] ), .S(n6386), .Y(n4883) );
  MUX2X1 U6062 ( .B(\Mem[42][10] ), .A(\Mem[43][10] ), .S(n6386), .Y(n4887) );
  MUX2X1 U6063 ( .B(\Mem[40][10] ), .A(\Mem[41][10] ), .S(n6386), .Y(n4886) );
  MUX2X1 U6064 ( .B(n4885), .A(n4882), .S(n6254), .Y(n4896) );
  MUX2X1 U6065 ( .B(\Mem[38][10] ), .A(\Mem[39][10] ), .S(n6386), .Y(n4890) );
  MUX2X1 U6066 ( .B(\Mem[36][10] ), .A(\Mem[37][10] ), .S(n6386), .Y(n4889) );
  MUX2X1 U6067 ( .B(\Mem[34][10] ), .A(\Mem[35][10] ), .S(n6386), .Y(n4893) );
  MUX2X1 U6068 ( .B(\Mem[32][10] ), .A(\Mem[33][10] ), .S(n6387), .Y(n4892) );
  MUX2X1 U6069 ( .B(n4891), .A(n4888), .S(n6254), .Y(n4895) );
  MUX2X1 U6070 ( .B(n4894), .A(n4879), .S(n6234), .Y(n4928) );
  MUX2X1 U6071 ( .B(\Mem[30][10] ), .A(\Mem[31][10] ), .S(n6387), .Y(n4899) );
  MUX2X1 U6072 ( .B(\Mem[28][10] ), .A(\Mem[29][10] ), .S(n6387), .Y(n4898) );
  MUX2X1 U6073 ( .B(\Mem[26][10] ), .A(\Mem[27][10] ), .S(n6387), .Y(n4902) );
  MUX2X1 U6074 ( .B(\Mem[24][10] ), .A(\Mem[25][10] ), .S(n6387), .Y(n4901) );
  MUX2X1 U6075 ( .B(n4900), .A(n4897), .S(n6254), .Y(n4911) );
  MUX2X1 U6076 ( .B(\Mem[22][10] ), .A(\Mem[23][10] ), .S(n6387), .Y(n4905) );
  MUX2X1 U6077 ( .B(\Mem[20][10] ), .A(\Mem[21][10] ), .S(n6387), .Y(n4904) );
  MUX2X1 U6078 ( .B(\Mem[18][10] ), .A(\Mem[19][10] ), .S(n6387), .Y(n4908) );
  MUX2X1 U6079 ( .B(\Mem[16][10] ), .A(\Mem[17][10] ), .S(n6387), .Y(n4907) );
  MUX2X1 U6080 ( .B(n4906), .A(n4903), .S(n6254), .Y(n4910) );
  MUX2X1 U6081 ( .B(\Mem[14][10] ), .A(\Mem[15][10] ), .S(n6387), .Y(n4914) );
  MUX2X1 U6082 ( .B(\Mem[12][10] ), .A(\Mem[13][10] ), .S(n6387), .Y(n4913) );
  MUX2X1 U6083 ( .B(\Mem[10][10] ), .A(\Mem[11][10] ), .S(n6387), .Y(n4917) );
  MUX2X1 U6084 ( .B(\Mem[8][10] ), .A(\Mem[9][10] ), .S(n6387), .Y(n4916) );
  MUX2X1 U6085 ( .B(n4915), .A(n4912), .S(n6254), .Y(n4926) );
  MUX2X1 U6086 ( .B(\Mem[6][10] ), .A(\Mem[7][10] ), .S(n6388), .Y(n4920) );
  MUX2X1 U6087 ( .B(\Mem[4][10] ), .A(\Mem[5][10] ), .S(n6388), .Y(n4919) );
  MUX2X1 U6088 ( .B(\Mem[2][10] ), .A(\Mem[3][10] ), .S(n6388), .Y(n4923) );
  MUX2X1 U6089 ( .B(\Mem[0][10] ), .A(\Mem[1][10] ), .S(n6388), .Y(n4922) );
  MUX2X1 U6090 ( .B(n4921), .A(n4918), .S(n6255), .Y(n4925) );
  MUX2X1 U6091 ( .B(n4924), .A(n4909), .S(n6234), .Y(n4927) );
  MUX2X1 U6092 ( .B(\Mem[62][11] ), .A(\Mem[63][11] ), .S(n6388), .Y(n4931) );
  MUX2X1 U6093 ( .B(\Mem[60][11] ), .A(\Mem[61][11] ), .S(n6388), .Y(n4930) );
  MUX2X1 U6094 ( .B(\Mem[58][11] ), .A(\Mem[59][11] ), .S(n6388), .Y(n4934) );
  MUX2X1 U6095 ( .B(\Mem[56][11] ), .A(\Mem[57][11] ), .S(n6388), .Y(n4933) );
  MUX2X1 U6096 ( .B(n4932), .A(n4929), .S(n6255), .Y(n4943) );
  MUX2X1 U6097 ( .B(\Mem[54][11] ), .A(\Mem[55][11] ), .S(n6388), .Y(n4937) );
  MUX2X1 U6098 ( .B(\Mem[52][11] ), .A(\Mem[53][11] ), .S(n6388), .Y(n4936) );
  MUX2X1 U6099 ( .B(\Mem[50][11] ), .A(\Mem[51][11] ), .S(n6388), .Y(n4940) );
  MUX2X1 U6100 ( .B(\Mem[48][11] ), .A(\Mem[49][11] ), .S(n6388), .Y(n4939) );
  MUX2X1 U6101 ( .B(n4938), .A(n4935), .S(n6255), .Y(n4942) );
  MUX2X1 U6102 ( .B(\Mem[46][11] ), .A(\Mem[47][11] ), .S(n6388), .Y(n4946) );
  MUX2X1 U6103 ( .B(\Mem[44][11] ), .A(\Mem[45][11] ), .S(n6389), .Y(n4945) );
  MUX2X1 U6104 ( .B(\Mem[42][11] ), .A(\Mem[43][11] ), .S(n6389), .Y(n4949) );
  MUX2X1 U6105 ( .B(\Mem[40][11] ), .A(\Mem[41][11] ), .S(n6389), .Y(n4948) );
  MUX2X1 U6106 ( .B(n4947), .A(n4944), .S(n6255), .Y(n4958) );
  MUX2X1 U6107 ( .B(\Mem[38][11] ), .A(\Mem[39][11] ), .S(n6389), .Y(n4952) );
  MUX2X1 U6108 ( .B(\Mem[36][11] ), .A(\Mem[37][11] ), .S(n6389), .Y(n4951) );
  MUX2X1 U6109 ( .B(\Mem[34][11] ), .A(\Mem[35][11] ), .S(n6389), .Y(n4955) );
  MUX2X1 U6110 ( .B(\Mem[32][11] ), .A(\Mem[33][11] ), .S(n6389), .Y(n4954) );
  MUX2X1 U6111 ( .B(n4953), .A(n4950), .S(n6255), .Y(n4957) );
  MUX2X1 U6112 ( .B(n4956), .A(n4941), .S(n6234), .Y(n4990) );
  MUX2X1 U6113 ( .B(\Mem[30][11] ), .A(\Mem[31][11] ), .S(n6389), .Y(n4961) );
  MUX2X1 U6114 ( .B(\Mem[28][11] ), .A(\Mem[29][11] ), .S(n6389), .Y(n4960) );
  MUX2X1 U6115 ( .B(\Mem[26][11] ), .A(\Mem[27][11] ), .S(n6389), .Y(n4964) );
  MUX2X1 U6116 ( .B(\Mem[24][11] ), .A(\Mem[25][11] ), .S(n6389), .Y(n4963) );
  MUX2X1 U6117 ( .B(n4962), .A(n4959), .S(n6255), .Y(n4973) );
  MUX2X1 U6118 ( .B(\Mem[22][11] ), .A(\Mem[23][11] ), .S(n6389), .Y(n4967) );
  MUX2X1 U6119 ( .B(\Mem[20][11] ), .A(\Mem[21][11] ), .S(n6389), .Y(n4966) );
  MUX2X1 U6120 ( .B(\Mem[18][11] ), .A(\Mem[19][11] ), .S(n6390), .Y(n4970) );
  MUX2X1 U6121 ( .B(\Mem[16][11] ), .A(\Mem[17][11] ), .S(n6390), .Y(n4969) );
  MUX2X1 U6122 ( .B(n4968), .A(n4965), .S(n6255), .Y(n4972) );
  MUX2X1 U6123 ( .B(\Mem[14][11] ), .A(\Mem[15][11] ), .S(n6390), .Y(n4976) );
  MUX2X1 U6124 ( .B(\Mem[12][11] ), .A(\Mem[13][11] ), .S(n6390), .Y(n4975) );
  MUX2X1 U6125 ( .B(\Mem[10][11] ), .A(\Mem[11][11] ), .S(n6390), .Y(n4979) );
  MUX2X1 U6126 ( .B(\Mem[8][11] ), .A(\Mem[9][11] ), .S(n6390), .Y(n4978) );
  MUX2X1 U6127 ( .B(n4977), .A(n4974), .S(n6255), .Y(n4988) );
  MUX2X1 U6128 ( .B(\Mem[6][11] ), .A(\Mem[7][11] ), .S(n6390), .Y(n4982) );
  MUX2X1 U6129 ( .B(\Mem[4][11] ), .A(\Mem[5][11] ), .S(n6390), .Y(n4981) );
  MUX2X1 U6130 ( .B(\Mem[2][11] ), .A(\Mem[3][11] ), .S(n6390), .Y(n4985) );
  MUX2X1 U6131 ( .B(\Mem[0][11] ), .A(\Mem[1][11] ), .S(n6390), .Y(n4984) );
  MUX2X1 U6132 ( .B(n4983), .A(n4980), .S(n6255), .Y(n4987) );
  MUX2X1 U6133 ( .B(n4986), .A(n4971), .S(n6234), .Y(n4989) );
  MUX2X1 U6134 ( .B(\Mem[62][12] ), .A(\Mem[63][12] ), .S(n6390), .Y(n4993) );
  MUX2X1 U6135 ( .B(\Mem[60][12] ), .A(\Mem[61][12] ), .S(n6390), .Y(n4992) );
  MUX2X1 U6136 ( .B(\Mem[58][12] ), .A(\Mem[59][12] ), .S(n6390), .Y(n4996) );
  MUX2X1 U6137 ( .B(\Mem[56][12] ), .A(\Mem[57][12] ), .S(n6391), .Y(n4995) );
  MUX2X1 U6138 ( .B(n4994), .A(n4991), .S(n6255), .Y(n5005) );
  MUX2X1 U6139 ( .B(\Mem[54][12] ), .A(\Mem[55][12] ), .S(n6391), .Y(n4999) );
  MUX2X1 U6140 ( .B(\Mem[52][12] ), .A(\Mem[53][12] ), .S(n6391), .Y(n4998) );
  MUX2X1 U6141 ( .B(\Mem[50][12] ), .A(\Mem[51][12] ), .S(n6391), .Y(n5002) );
  MUX2X1 U6142 ( .B(\Mem[48][12] ), .A(\Mem[49][12] ), .S(n6391), .Y(n5001) );
  MUX2X1 U6143 ( .B(n5000), .A(n4997), .S(n6255), .Y(n5004) );
  MUX2X1 U6144 ( .B(\Mem[46][12] ), .A(\Mem[47][12] ), .S(n6391), .Y(n5008) );
  MUX2X1 U6145 ( .B(\Mem[44][12] ), .A(\Mem[45][12] ), .S(n6391), .Y(n5007) );
  MUX2X1 U6146 ( .B(\Mem[42][12] ), .A(\Mem[43][12] ), .S(n6391), .Y(n5011) );
  MUX2X1 U6147 ( .B(\Mem[40][12] ), .A(\Mem[41][12] ), .S(n6391), .Y(n5010) );
  MUX2X1 U6148 ( .B(n5009), .A(n5006), .S(n6255), .Y(n5020) );
  MUX2X1 U6149 ( .B(\Mem[38][12] ), .A(\Mem[39][12] ), .S(n6391), .Y(n5014) );
  MUX2X1 U6150 ( .B(\Mem[36][12] ), .A(\Mem[37][12] ), .S(n6391), .Y(n5013) );
  MUX2X1 U6151 ( .B(\Mem[34][12] ), .A(\Mem[35][12] ), .S(n6391), .Y(n5017) );
  MUX2X1 U6152 ( .B(\Mem[32][12] ), .A(\Mem[33][12] ), .S(n6391), .Y(n5016) );
  MUX2X1 U6153 ( .B(n5015), .A(n5012), .S(n6255), .Y(n5019) );
  MUX2X1 U6154 ( .B(n5018), .A(n5003), .S(n6234), .Y(n5052) );
  MUX2X1 U6155 ( .B(\Mem[30][12] ), .A(\Mem[31][12] ), .S(n6392), .Y(n5023) );
  MUX2X1 U6156 ( .B(\Mem[28][12] ), .A(\Mem[29][12] ), .S(n6392), .Y(n5022) );
  MUX2X1 U6157 ( .B(\Mem[26][12] ), .A(\Mem[27][12] ), .S(n6392), .Y(n5026) );
  MUX2X1 U6158 ( .B(\Mem[24][12] ), .A(\Mem[25][12] ), .S(n6392), .Y(n5025) );
  MUX2X1 U6159 ( .B(n5024), .A(n5021), .S(n6256), .Y(n5035) );
  MUX2X1 U6160 ( .B(\Mem[22][12] ), .A(\Mem[23][12] ), .S(n6392), .Y(n5029) );
  MUX2X1 U6161 ( .B(\Mem[20][12] ), .A(\Mem[21][12] ), .S(n6392), .Y(n5028) );
  MUX2X1 U6162 ( .B(\Mem[18][12] ), .A(\Mem[19][12] ), .S(n6392), .Y(n5032) );
  MUX2X1 U6163 ( .B(\Mem[16][12] ), .A(\Mem[17][12] ), .S(n6392), .Y(n5031) );
  MUX2X1 U6164 ( .B(n5030), .A(n5027), .S(n6256), .Y(n5034) );
  MUX2X1 U6165 ( .B(\Mem[14][12] ), .A(\Mem[15][12] ), .S(n6392), .Y(n5038) );
  MUX2X1 U6166 ( .B(\Mem[12][12] ), .A(\Mem[13][12] ), .S(n6392), .Y(n5037) );
  MUX2X1 U6167 ( .B(\Mem[10][12] ), .A(\Mem[11][12] ), .S(n6392), .Y(n5041) );
  MUX2X1 U6168 ( .B(\Mem[8][12] ), .A(\Mem[9][12] ), .S(n6392), .Y(n5040) );
  MUX2X1 U6169 ( .B(n5039), .A(n5036), .S(n6256), .Y(n5050) );
  MUX2X1 U6170 ( .B(\Mem[6][12] ), .A(\Mem[7][12] ), .S(n6392), .Y(n5044) );
  MUX2X1 U6171 ( .B(\Mem[4][12] ), .A(\Mem[5][12] ), .S(n6393), .Y(n5043) );
  MUX2X1 U6172 ( .B(\Mem[2][12] ), .A(\Mem[3][12] ), .S(n6393), .Y(n5047) );
  MUX2X1 U6173 ( .B(\Mem[0][12] ), .A(\Mem[1][12] ), .S(n6393), .Y(n5046) );
  MUX2X1 U6174 ( .B(n5045), .A(n5042), .S(n6256), .Y(n5049) );
  MUX2X1 U6175 ( .B(n5048), .A(n5033), .S(n6235), .Y(n5051) );
  MUX2X1 U6176 ( .B(\Mem[62][13] ), .A(\Mem[63][13] ), .S(n6393), .Y(n5055) );
  MUX2X1 U6177 ( .B(\Mem[60][13] ), .A(\Mem[61][13] ), .S(n6393), .Y(n5054) );
  MUX2X1 U6178 ( .B(\Mem[58][13] ), .A(\Mem[59][13] ), .S(n6393), .Y(n5058) );
  MUX2X1 U6179 ( .B(\Mem[56][13] ), .A(\Mem[57][13] ), .S(n6393), .Y(n5057) );
  MUX2X1 U6180 ( .B(n5056), .A(n5053), .S(n6256), .Y(n5067) );
  MUX2X1 U6181 ( .B(\Mem[54][13] ), .A(\Mem[55][13] ), .S(n6393), .Y(n5061) );
  MUX2X1 U6182 ( .B(\Mem[52][13] ), .A(\Mem[53][13] ), .S(n6393), .Y(n5060) );
  MUX2X1 U6183 ( .B(\Mem[50][13] ), .A(\Mem[51][13] ), .S(n6393), .Y(n5064) );
  MUX2X1 U6184 ( .B(\Mem[48][13] ), .A(\Mem[49][13] ), .S(n6393), .Y(n5063) );
  MUX2X1 U6185 ( .B(n5062), .A(n5059), .S(n6256), .Y(n5066) );
  MUX2X1 U6186 ( .B(\Mem[46][13] ), .A(\Mem[47][13] ), .S(n6393), .Y(n5070) );
  MUX2X1 U6187 ( .B(\Mem[44][13] ), .A(\Mem[45][13] ), .S(n6393), .Y(n5069) );
  MUX2X1 U6188 ( .B(\Mem[42][13] ), .A(\Mem[43][13] ), .S(n6394), .Y(n5073) );
  MUX2X1 U6189 ( .B(\Mem[40][13] ), .A(\Mem[41][13] ), .S(n6394), .Y(n5072) );
  MUX2X1 U6190 ( .B(n5071), .A(n5068), .S(n6256), .Y(n5082) );
  MUX2X1 U6191 ( .B(\Mem[38][13] ), .A(\Mem[39][13] ), .S(n6394), .Y(n5076) );
  MUX2X1 U6192 ( .B(\Mem[36][13] ), .A(\Mem[37][13] ), .S(n6394), .Y(n5075) );
  MUX2X1 U6193 ( .B(\Mem[34][13] ), .A(\Mem[35][13] ), .S(n6394), .Y(n5079) );
  MUX2X1 U6194 ( .B(\Mem[32][13] ), .A(\Mem[33][13] ), .S(n6394), .Y(n5078) );
  MUX2X1 U6195 ( .B(n5077), .A(n5074), .S(n6256), .Y(n5081) );
  MUX2X1 U6196 ( .B(n5080), .A(n5065), .S(n6235), .Y(n5114) );
  MUX2X1 U6197 ( .B(\Mem[30][13] ), .A(\Mem[31][13] ), .S(n6394), .Y(n5085) );
  MUX2X1 U6198 ( .B(\Mem[28][13] ), .A(\Mem[29][13] ), .S(n6394), .Y(n5084) );
  MUX2X1 U6199 ( .B(\Mem[26][13] ), .A(\Mem[27][13] ), .S(n6394), .Y(n5088) );
  MUX2X1 U6200 ( .B(\Mem[24][13] ), .A(\Mem[25][13] ), .S(n6394), .Y(n5087) );
  MUX2X1 U6201 ( .B(n5086), .A(n5083), .S(n6256), .Y(n5097) );
  MUX2X1 U6202 ( .B(\Mem[22][13] ), .A(\Mem[23][13] ), .S(n6394), .Y(n5091) );
  MUX2X1 U6203 ( .B(\Mem[20][13] ), .A(\Mem[21][13] ), .S(n6394), .Y(n5090) );
  MUX2X1 U6204 ( .B(\Mem[18][13] ), .A(\Mem[19][13] ), .S(n6394), .Y(n5094) );
  MUX2X1 U6205 ( .B(\Mem[16][13] ), .A(\Mem[17][13] ), .S(n6395), .Y(n5093) );
  MUX2X1 U6206 ( .B(n5092), .A(n5089), .S(n6256), .Y(n5096) );
  MUX2X1 U6207 ( .B(\Mem[14][13] ), .A(\Mem[15][13] ), .S(n6395), .Y(n5100) );
  MUX2X1 U6208 ( .B(\Mem[12][13] ), .A(\Mem[13][13] ), .S(n6395), .Y(n5099) );
  MUX2X1 U6209 ( .B(\Mem[10][13] ), .A(\Mem[11][13] ), .S(n6395), .Y(n5103) );
  MUX2X1 U6210 ( .B(\Mem[8][13] ), .A(\Mem[9][13] ), .S(n6395), .Y(n5102) );
  MUX2X1 U6211 ( .B(n5101), .A(n5098), .S(n6256), .Y(n5112) );
  MUX2X1 U6212 ( .B(\Mem[6][13] ), .A(\Mem[7][13] ), .S(n6395), .Y(n5106) );
  MUX2X1 U6213 ( .B(\Mem[4][13] ), .A(\Mem[5][13] ), .S(n6395), .Y(n5105) );
  MUX2X1 U6214 ( .B(\Mem[2][13] ), .A(\Mem[3][13] ), .S(n6395), .Y(n5109) );
  MUX2X1 U6215 ( .B(\Mem[0][13] ), .A(\Mem[1][13] ), .S(n6395), .Y(n5108) );
  MUX2X1 U6216 ( .B(n5107), .A(n5104), .S(n6256), .Y(n5111) );
  MUX2X1 U6217 ( .B(n5110), .A(n5095), .S(n6235), .Y(n5113) );
  MUX2X1 U6218 ( .B(\Mem[62][14] ), .A(\Mem[63][14] ), .S(n6395), .Y(n5117) );
  MUX2X1 U6219 ( .B(\Mem[60][14] ), .A(\Mem[61][14] ), .S(n6395), .Y(n5116) );
  MUX2X1 U6220 ( .B(\Mem[58][14] ), .A(\Mem[59][14] ), .S(n6395), .Y(n5120) );
  MUX2X1 U6221 ( .B(\Mem[56][14] ), .A(\Mem[57][14] ), .S(n6395), .Y(n5119) );
  MUX2X1 U6222 ( .B(n5118), .A(n5115), .S(n6256), .Y(n5129) );
  MUX2X1 U6223 ( .B(\Mem[54][14] ), .A(\Mem[55][14] ), .S(n6396), .Y(n5123) );
  MUX2X1 U6224 ( .B(\Mem[52][14] ), .A(\Mem[53][14] ), .S(n6396), .Y(n5122) );
  MUX2X1 U6225 ( .B(\Mem[50][14] ), .A(\Mem[51][14] ), .S(n6396), .Y(n5126) );
  MUX2X1 U6226 ( .B(\Mem[48][14] ), .A(\Mem[49][14] ), .S(n6396), .Y(n5125) );
  MUX2X1 U6227 ( .B(n5124), .A(n5121), .S(n6257), .Y(n5128) );
  MUX2X1 U6228 ( .B(\Mem[46][14] ), .A(\Mem[47][14] ), .S(n6396), .Y(n5132) );
  MUX2X1 U6229 ( .B(\Mem[44][14] ), .A(\Mem[45][14] ), .S(n6396), .Y(n5131) );
  MUX2X1 U6230 ( .B(\Mem[42][14] ), .A(\Mem[43][14] ), .S(n6396), .Y(n5135) );
  MUX2X1 U6231 ( .B(\Mem[40][14] ), .A(\Mem[41][14] ), .S(n6396), .Y(n5134) );
  MUX2X1 U6232 ( .B(n5133), .A(n5130), .S(n6257), .Y(n5144) );
  MUX2X1 U6233 ( .B(\Mem[38][14] ), .A(\Mem[39][14] ), .S(n6396), .Y(n5138) );
  MUX2X1 U6234 ( .B(\Mem[36][14] ), .A(\Mem[37][14] ), .S(n6396), .Y(n5137) );
  MUX2X1 U6235 ( .B(\Mem[34][14] ), .A(\Mem[35][14] ), .S(n6396), .Y(n5141) );
  MUX2X1 U6236 ( .B(\Mem[32][14] ), .A(\Mem[33][14] ), .S(n6396), .Y(n5140) );
  MUX2X1 U6237 ( .B(n5139), .A(n5136), .S(n6257), .Y(n5143) );
  MUX2X1 U6238 ( .B(n5142), .A(n5127), .S(n6235), .Y(n5176) );
  MUX2X1 U6239 ( .B(\Mem[30][14] ), .A(\Mem[31][14] ), .S(n6396), .Y(n5147) );
  MUX2X1 U6240 ( .B(\Mem[28][14] ), .A(\Mem[29][14] ), .S(n6397), .Y(n5146) );
  MUX2X1 U6241 ( .B(\Mem[26][14] ), .A(\Mem[27][14] ), .S(n6397), .Y(n5150) );
  MUX2X1 U6242 ( .B(\Mem[24][14] ), .A(\Mem[25][14] ), .S(n6397), .Y(n5149) );
  MUX2X1 U6243 ( .B(n5148), .A(n5145), .S(n6257), .Y(n5159) );
  MUX2X1 U6244 ( .B(\Mem[22][14] ), .A(\Mem[23][14] ), .S(n6397), .Y(n5153) );
  MUX2X1 U6245 ( .B(\Mem[20][14] ), .A(\Mem[21][14] ), .S(n6397), .Y(n5152) );
  MUX2X1 U6246 ( .B(\Mem[18][14] ), .A(\Mem[19][14] ), .S(n6397), .Y(n5156) );
  MUX2X1 U6247 ( .B(\Mem[16][14] ), .A(\Mem[17][14] ), .S(n6397), .Y(n5155) );
  MUX2X1 U6248 ( .B(n5154), .A(n5151), .S(n6257), .Y(n5158) );
  MUX2X1 U6249 ( .B(\Mem[14][14] ), .A(\Mem[15][14] ), .S(n6397), .Y(n5162) );
  MUX2X1 U6250 ( .B(\Mem[12][14] ), .A(\Mem[13][14] ), .S(n6397), .Y(n5161) );
  MUX2X1 U6251 ( .B(\Mem[10][14] ), .A(\Mem[11][14] ), .S(n6397), .Y(n5165) );
  MUX2X1 U6252 ( .B(\Mem[8][14] ), .A(\Mem[9][14] ), .S(n6397), .Y(n5164) );
  MUX2X1 U6253 ( .B(n5163), .A(n5160), .S(n6257), .Y(n5174) );
  MUX2X1 U6254 ( .B(\Mem[6][14] ), .A(\Mem[7][14] ), .S(n6397), .Y(n5168) );
  MUX2X1 U6255 ( .B(\Mem[4][14] ), .A(\Mem[5][14] ), .S(n6397), .Y(n5167) );
  MUX2X1 U6256 ( .B(\Mem[2][14] ), .A(\Mem[3][14] ), .S(n6398), .Y(n5171) );
  MUX2X1 U6257 ( .B(\Mem[0][14] ), .A(\Mem[1][14] ), .S(n6398), .Y(n5170) );
  MUX2X1 U6258 ( .B(n5169), .A(n5166), .S(n6257), .Y(n5173) );
  MUX2X1 U6259 ( .B(n5172), .A(n5157), .S(n6235), .Y(n5175) );
  MUX2X1 U6260 ( .B(\Mem[62][15] ), .A(\Mem[63][15] ), .S(n6398), .Y(n5179) );
  MUX2X1 U6261 ( .B(\Mem[60][15] ), .A(\Mem[61][15] ), .S(n6398), .Y(n5178) );
  MUX2X1 U6262 ( .B(\Mem[58][15] ), .A(\Mem[59][15] ), .S(n6398), .Y(n5182) );
  MUX2X1 U6263 ( .B(\Mem[56][15] ), .A(\Mem[57][15] ), .S(n6398), .Y(n5181) );
  MUX2X1 U6264 ( .B(n5180), .A(n5177), .S(n6257), .Y(n5191) );
  MUX2X1 U6265 ( .B(\Mem[54][15] ), .A(\Mem[55][15] ), .S(n6398), .Y(n5185) );
  MUX2X1 U6266 ( .B(\Mem[52][15] ), .A(\Mem[53][15] ), .S(n6398), .Y(n5184) );
  MUX2X1 U6267 ( .B(\Mem[50][15] ), .A(\Mem[51][15] ), .S(n6398), .Y(n5188) );
  MUX2X1 U6268 ( .B(\Mem[48][15] ), .A(\Mem[49][15] ), .S(n6398), .Y(n5187) );
  MUX2X1 U6269 ( .B(n5186), .A(n5183), .S(n6257), .Y(n5190) );
  MUX2X1 U6270 ( .B(\Mem[46][15] ), .A(\Mem[47][15] ), .S(n6398), .Y(n5194) );
  MUX2X1 U6271 ( .B(\Mem[44][15] ), .A(\Mem[45][15] ), .S(n6398), .Y(n5193) );
  MUX2X1 U6272 ( .B(\Mem[42][15] ), .A(\Mem[43][15] ), .S(n6398), .Y(n5197) );
  MUX2X1 U6273 ( .B(\Mem[40][15] ), .A(\Mem[41][15] ), .S(n6399), .Y(n5196) );
  MUX2X1 U6274 ( .B(n5195), .A(n5192), .S(n6257), .Y(n5206) );
  MUX2X1 U6275 ( .B(\Mem[38][15] ), .A(\Mem[39][15] ), .S(n6399), .Y(n5200) );
  MUX2X1 U6276 ( .B(\Mem[36][15] ), .A(\Mem[37][15] ), .S(n6399), .Y(n5199) );
  MUX2X1 U6277 ( .B(\Mem[34][15] ), .A(\Mem[35][15] ), .S(n6399), .Y(n5203) );
  MUX2X1 U6278 ( .B(\Mem[32][15] ), .A(\Mem[33][15] ), .S(n6399), .Y(n5202) );
  MUX2X1 U6279 ( .B(n5201), .A(n5198), .S(n6257), .Y(n5205) );
  MUX2X1 U6280 ( .B(n5204), .A(n5189), .S(n6235), .Y(n5238) );
  MUX2X1 U6281 ( .B(\Mem[30][15] ), .A(\Mem[31][15] ), .S(n6399), .Y(n5209) );
  MUX2X1 U6282 ( .B(\Mem[28][15] ), .A(\Mem[29][15] ), .S(n6399), .Y(n5208) );
  MUX2X1 U6283 ( .B(\Mem[26][15] ), .A(\Mem[27][15] ), .S(n6399), .Y(n5212) );
  MUX2X1 U6284 ( .B(\Mem[24][15] ), .A(\Mem[25][15] ), .S(n6399), .Y(n5211) );
  MUX2X1 U6285 ( .B(n5210), .A(n5207), .S(n6257), .Y(n5221) );
  MUX2X1 U6286 ( .B(\Mem[22][15] ), .A(\Mem[23][15] ), .S(n6399), .Y(n5215) );
  MUX2X1 U6287 ( .B(\Mem[20][15] ), .A(\Mem[21][15] ), .S(n6399), .Y(n5214) );
  MUX2X1 U6288 ( .B(\Mem[18][15] ), .A(\Mem[19][15] ), .S(n6399), .Y(n5218) );
  MUX2X1 U6289 ( .B(\Mem[16][15] ), .A(\Mem[17][15] ), .S(n6399), .Y(n5217) );
  MUX2X1 U6290 ( .B(n5216), .A(n5213), .S(n6257), .Y(n5220) );
  MUX2X1 U6291 ( .B(\Mem[14][15] ), .A(\Mem[15][15] ), .S(n6400), .Y(n5224) );
  MUX2X1 U6292 ( .B(\Mem[12][15] ), .A(\Mem[13][15] ), .S(n6400), .Y(n5223) );
  MUX2X1 U6293 ( .B(\Mem[10][15] ), .A(\Mem[11][15] ), .S(n6400), .Y(n5227) );
  MUX2X1 U6294 ( .B(\Mem[8][15] ), .A(\Mem[9][15] ), .S(n6400), .Y(n5226) );
  MUX2X1 U6295 ( .B(n5225), .A(n5222), .S(n6258), .Y(n5236) );
  MUX2X1 U6296 ( .B(\Mem[6][15] ), .A(\Mem[7][15] ), .S(n6400), .Y(n5230) );
  MUX2X1 U6297 ( .B(\Mem[4][15] ), .A(\Mem[5][15] ), .S(n6400), .Y(n5229) );
  MUX2X1 U6298 ( .B(\Mem[2][15] ), .A(\Mem[3][15] ), .S(n6400), .Y(n5233) );
  MUX2X1 U6299 ( .B(\Mem[0][15] ), .A(\Mem[1][15] ), .S(n6400), .Y(n5232) );
  MUX2X1 U6300 ( .B(n5231), .A(n5228), .S(n6258), .Y(n5235) );
  MUX2X1 U6301 ( .B(n5234), .A(n5219), .S(n6235), .Y(n5237) );
  MUX2X1 U6302 ( .B(\Mem[62][16] ), .A(\Mem[63][16] ), .S(n6400), .Y(n5241) );
  MUX2X1 U6303 ( .B(\Mem[60][16] ), .A(\Mem[61][16] ), .S(n6400), .Y(n5240) );
  MUX2X1 U6304 ( .B(\Mem[58][16] ), .A(\Mem[59][16] ), .S(n6400), .Y(n5244) );
  MUX2X1 U6305 ( .B(\Mem[56][16] ), .A(\Mem[57][16] ), .S(n6400), .Y(n5243) );
  MUX2X1 U6306 ( .B(n5242), .A(n5239), .S(n6258), .Y(n5253) );
  MUX2X1 U6307 ( .B(\Mem[54][16] ), .A(\Mem[55][16] ), .S(n6400), .Y(n5247) );
  MUX2X1 U6308 ( .B(\Mem[52][16] ), .A(\Mem[53][16] ), .S(n6401), .Y(n5246) );
  MUX2X1 U6309 ( .B(\Mem[50][16] ), .A(\Mem[51][16] ), .S(n6401), .Y(n5250) );
  MUX2X1 U6310 ( .B(\Mem[48][16] ), .A(\Mem[49][16] ), .S(n6401), .Y(n5249) );
  MUX2X1 U6311 ( .B(n5248), .A(n5245), .S(n6258), .Y(n5252) );
  MUX2X1 U6312 ( .B(\Mem[46][16] ), .A(\Mem[47][16] ), .S(n6401), .Y(n5256) );
  MUX2X1 U6313 ( .B(\Mem[44][16] ), .A(\Mem[45][16] ), .S(n6401), .Y(n5255) );
  MUX2X1 U6314 ( .B(\Mem[42][16] ), .A(\Mem[43][16] ), .S(n6401), .Y(n5259) );
  MUX2X1 U6315 ( .B(\Mem[40][16] ), .A(\Mem[41][16] ), .S(n6401), .Y(n5258) );
  MUX2X1 U6316 ( .B(n5257), .A(n5254), .S(n6258), .Y(n5268) );
  MUX2X1 U6317 ( .B(\Mem[38][16] ), .A(\Mem[39][16] ), .S(n6401), .Y(n5262) );
  MUX2X1 U6318 ( .B(\Mem[36][16] ), .A(\Mem[37][16] ), .S(n6401), .Y(n5261) );
  MUX2X1 U6319 ( .B(\Mem[34][16] ), .A(\Mem[35][16] ), .S(n6401), .Y(n5265) );
  MUX2X1 U6320 ( .B(\Mem[32][16] ), .A(\Mem[33][16] ), .S(n6401), .Y(n5264) );
  MUX2X1 U6321 ( .B(n5263), .A(n5260), .S(n6258), .Y(n5267) );
  MUX2X1 U6322 ( .B(n5266), .A(n5251), .S(n6235), .Y(n5300) );
  MUX2X1 U6323 ( .B(\Mem[30][16] ), .A(\Mem[31][16] ), .S(n6401), .Y(n5271) );
  MUX2X1 U6324 ( .B(\Mem[28][16] ), .A(\Mem[29][16] ), .S(n6401), .Y(n5270) );
  MUX2X1 U6325 ( .B(\Mem[26][16] ), .A(\Mem[27][16] ), .S(n6402), .Y(n5274) );
  MUX2X1 U6326 ( .B(\Mem[24][16] ), .A(\Mem[25][16] ), .S(n6402), .Y(n5273) );
  MUX2X1 U6327 ( .B(n5272), .A(n5269), .S(n6258), .Y(n5283) );
  MUX2X1 U6328 ( .B(\Mem[22][16] ), .A(\Mem[23][16] ), .S(n6402), .Y(n5277) );
  MUX2X1 U6329 ( .B(\Mem[20][16] ), .A(\Mem[21][16] ), .S(n6402), .Y(n5276) );
  MUX2X1 U6330 ( .B(\Mem[18][16] ), .A(\Mem[19][16] ), .S(n6402), .Y(n5280) );
  MUX2X1 U6331 ( .B(\Mem[16][16] ), .A(\Mem[17][16] ), .S(n6402), .Y(n5279) );
  MUX2X1 U6332 ( .B(n5278), .A(n5275), .S(n6258), .Y(n5282) );
  MUX2X1 U6333 ( .B(\Mem[14][16] ), .A(\Mem[15][16] ), .S(n6402), .Y(n5286) );
  MUX2X1 U6334 ( .B(\Mem[12][16] ), .A(\Mem[13][16] ), .S(n6402), .Y(n5285) );
  MUX2X1 U6335 ( .B(\Mem[10][16] ), .A(\Mem[11][16] ), .S(n6402), .Y(n5289) );
  MUX2X1 U6336 ( .B(\Mem[8][16] ), .A(\Mem[9][16] ), .S(n6402), .Y(n5288) );
  MUX2X1 U6337 ( .B(n5287), .A(n5284), .S(n6258), .Y(n5298) );
  MUX2X1 U6338 ( .B(\Mem[6][16] ), .A(\Mem[7][16] ), .S(n6402), .Y(n5292) );
  MUX2X1 U6339 ( .B(\Mem[4][16] ), .A(\Mem[5][16] ), .S(n6402), .Y(n5291) );
  MUX2X1 U6340 ( .B(\Mem[2][16] ), .A(\Mem[3][16] ), .S(n6402), .Y(n5295) );
  MUX2X1 U6341 ( .B(\Mem[0][16] ), .A(\Mem[1][16] ), .S(n6403), .Y(n5294) );
  MUX2X1 U6342 ( .B(n5293), .A(n5290), .S(n6258), .Y(n5297) );
  MUX2X1 U6343 ( .B(n5296), .A(n5281), .S(n6235), .Y(n5299) );
  MUX2X1 U6344 ( .B(\Mem[62][17] ), .A(\Mem[63][17] ), .S(n6403), .Y(n5303) );
  MUX2X1 U6345 ( .B(\Mem[60][17] ), .A(\Mem[61][17] ), .S(n6403), .Y(n5302) );
  MUX2X1 U6346 ( .B(\Mem[58][17] ), .A(\Mem[59][17] ), .S(n6403), .Y(n5306) );
  MUX2X1 U6347 ( .B(\Mem[56][17] ), .A(\Mem[57][17] ), .S(n6403), .Y(n5305) );
  MUX2X1 U6348 ( .B(n5304), .A(n5301), .S(n6258), .Y(n5315) );
  MUX2X1 U6349 ( .B(\Mem[54][17] ), .A(\Mem[55][17] ), .S(n6403), .Y(n5309) );
  MUX2X1 U6350 ( .B(\Mem[52][17] ), .A(\Mem[53][17] ), .S(n6403), .Y(n5308) );
  MUX2X1 U6351 ( .B(\Mem[50][17] ), .A(\Mem[51][17] ), .S(n6403), .Y(n5312) );
  MUX2X1 U6352 ( .B(\Mem[48][17] ), .A(\Mem[49][17] ), .S(n6403), .Y(n5311) );
  MUX2X1 U6353 ( .B(n5310), .A(n5307), .S(n6258), .Y(n5314) );
  MUX2X1 U6354 ( .B(\Mem[46][17] ), .A(\Mem[47][17] ), .S(n6403), .Y(n5318) );
  MUX2X1 U6355 ( .B(\Mem[44][17] ), .A(\Mem[45][17] ), .S(n6403), .Y(n5317) );
  MUX2X1 U6356 ( .B(\Mem[42][17] ), .A(\Mem[43][17] ), .S(n6403), .Y(n5321) );
  MUX2X1 U6357 ( .B(\Mem[40][17] ), .A(\Mem[41][17] ), .S(n6403), .Y(n5320) );
  MUX2X1 U6358 ( .B(n5319), .A(n5316), .S(n6258), .Y(n5330) );
  MUX2X1 U6359 ( .B(\Mem[38][17] ), .A(\Mem[39][17] ), .S(n6404), .Y(n5324) );
  MUX2X1 U6360 ( .B(\Mem[36][17] ), .A(\Mem[37][17] ), .S(n6404), .Y(n5323) );
  MUX2X1 U6361 ( .B(\Mem[34][17] ), .A(\Mem[35][17] ), .S(n6404), .Y(n5327) );
  MUX2X1 U6362 ( .B(\Mem[32][17] ), .A(\Mem[33][17] ), .S(n6404), .Y(n5326) );
  MUX2X1 U6363 ( .B(n5325), .A(n5322), .S(n6259), .Y(n5329) );
  MUX2X1 U6364 ( .B(n5328), .A(n5313), .S(n6235), .Y(n5362) );
  MUX2X1 U6365 ( .B(\Mem[30][17] ), .A(\Mem[31][17] ), .S(n6404), .Y(n5333) );
  MUX2X1 U6366 ( .B(\Mem[28][17] ), .A(\Mem[29][17] ), .S(n6404), .Y(n5332) );
  MUX2X1 U6367 ( .B(\Mem[26][17] ), .A(\Mem[27][17] ), .S(n6404), .Y(n5336) );
  MUX2X1 U6368 ( .B(\Mem[24][17] ), .A(\Mem[25][17] ), .S(n6404), .Y(n5335) );
  MUX2X1 U6369 ( .B(n5334), .A(n5331), .S(n6259), .Y(n5345) );
  MUX2X1 U6370 ( .B(\Mem[22][17] ), .A(\Mem[23][17] ), .S(n6404), .Y(n5339) );
  MUX2X1 U6371 ( .B(\Mem[20][17] ), .A(\Mem[21][17] ), .S(n6404), .Y(n5338) );
  MUX2X1 U6372 ( .B(\Mem[18][17] ), .A(\Mem[19][17] ), .S(n6404), .Y(n5342) );
  MUX2X1 U6373 ( .B(\Mem[16][17] ), .A(\Mem[17][17] ), .S(n6404), .Y(n5341) );
  MUX2X1 U6374 ( .B(n5340), .A(n5337), .S(n6259), .Y(n5344) );
  MUX2X1 U6375 ( .B(\Mem[14][17] ), .A(\Mem[15][17] ), .S(n6404), .Y(n5348) );
  MUX2X1 U6376 ( .B(\Mem[12][17] ), .A(\Mem[13][17] ), .S(n6405), .Y(n5347) );
  MUX2X1 U6377 ( .B(\Mem[10][17] ), .A(\Mem[11][17] ), .S(n6405), .Y(n5351) );
  MUX2X1 U6378 ( .B(\Mem[8][17] ), .A(\Mem[9][17] ), .S(n6405), .Y(n5350) );
  MUX2X1 U6379 ( .B(n5349), .A(n5346), .S(n6259), .Y(n5360) );
  MUX2X1 U6380 ( .B(\Mem[6][17] ), .A(\Mem[7][17] ), .S(n6405), .Y(n5354) );
  MUX2X1 U6381 ( .B(\Mem[4][17] ), .A(\Mem[5][17] ), .S(n6405), .Y(n5353) );
  MUX2X1 U6382 ( .B(\Mem[2][17] ), .A(\Mem[3][17] ), .S(n6405), .Y(n5357) );
  MUX2X1 U6383 ( .B(\Mem[0][17] ), .A(\Mem[1][17] ), .S(n6405), .Y(n5356) );
  MUX2X1 U6384 ( .B(n5355), .A(n5352), .S(n6259), .Y(n5359) );
  MUX2X1 U6385 ( .B(n5358), .A(n5343), .S(n6235), .Y(n5361) );
  MUX2X1 U6386 ( .B(\Mem[62][18] ), .A(\Mem[63][18] ), .S(n6405), .Y(n5365) );
  MUX2X1 U6387 ( .B(\Mem[60][18] ), .A(\Mem[61][18] ), .S(n6405), .Y(n5364) );
  MUX2X1 U6388 ( .B(\Mem[58][18] ), .A(\Mem[59][18] ), .S(n6405), .Y(n5368) );
  MUX2X1 U6389 ( .B(\Mem[56][18] ), .A(\Mem[57][18] ), .S(n6405), .Y(n5367) );
  MUX2X1 U6390 ( .B(n5366), .A(n5363), .S(n6259), .Y(n5377) );
  MUX2X1 U6391 ( .B(\Mem[54][18] ), .A(\Mem[55][18] ), .S(n6405), .Y(n5371) );
  MUX2X1 U6392 ( .B(\Mem[52][18] ), .A(\Mem[53][18] ), .S(n6405), .Y(n5370) );
  MUX2X1 U6393 ( .B(\Mem[50][18] ), .A(\Mem[51][18] ), .S(n6406), .Y(n5374) );
  MUX2X1 U6394 ( .B(\Mem[48][18] ), .A(\Mem[49][18] ), .S(n6406), .Y(n5373) );
  MUX2X1 U6395 ( .B(n5372), .A(n5369), .S(n6259), .Y(n5376) );
  MUX2X1 U6396 ( .B(\Mem[46][18] ), .A(\Mem[47][18] ), .S(n6406), .Y(n5380) );
  MUX2X1 U6397 ( .B(\Mem[44][18] ), .A(\Mem[45][18] ), .S(n6406), .Y(n5379) );
  MUX2X1 U6398 ( .B(\Mem[42][18] ), .A(\Mem[43][18] ), .S(n6406), .Y(n5383) );
  MUX2X1 U6399 ( .B(\Mem[40][18] ), .A(\Mem[41][18] ), .S(n6406), .Y(n5382) );
  MUX2X1 U6400 ( .B(n5381), .A(n5378), .S(n6259), .Y(n5392) );
  MUX2X1 U6401 ( .B(\Mem[38][18] ), .A(\Mem[39][18] ), .S(n6406), .Y(n5386) );
  MUX2X1 U6402 ( .B(\Mem[36][18] ), .A(\Mem[37][18] ), .S(n6406), .Y(n5385) );
  MUX2X1 U6403 ( .B(\Mem[34][18] ), .A(\Mem[35][18] ), .S(n6406), .Y(n5389) );
  MUX2X1 U6404 ( .B(\Mem[32][18] ), .A(\Mem[33][18] ), .S(n6406), .Y(n5388) );
  MUX2X1 U6405 ( .B(n5387), .A(n5384), .S(n6259), .Y(n5391) );
  MUX2X1 U6406 ( .B(n5390), .A(n5375), .S(n6235), .Y(n5424) );
  MUX2X1 U6407 ( .B(\Mem[30][18] ), .A(\Mem[31][18] ), .S(n6406), .Y(n5395) );
  MUX2X1 U6408 ( .B(\Mem[28][18] ), .A(\Mem[29][18] ), .S(n6406), .Y(n5394) );
  MUX2X1 U6409 ( .B(\Mem[26][18] ), .A(\Mem[27][18] ), .S(n6406), .Y(n5398) );
  MUX2X1 U6410 ( .B(\Mem[24][18] ), .A(\Mem[25][18] ), .S(n6407), .Y(n5397) );
  MUX2X1 U6411 ( .B(n5396), .A(n5393), .S(n6259), .Y(n5407) );
  MUX2X1 U6412 ( .B(\Mem[22][18] ), .A(\Mem[23][18] ), .S(n6407), .Y(n5401) );
  MUX2X1 U6413 ( .B(\Mem[20][18] ), .A(\Mem[21][18] ), .S(n6407), .Y(n5400) );
  MUX2X1 U6414 ( .B(\Mem[18][18] ), .A(\Mem[19][18] ), .S(n6407), .Y(n5404) );
  MUX2X1 U6415 ( .B(\Mem[16][18] ), .A(\Mem[17][18] ), .S(n6407), .Y(n5403) );
  MUX2X1 U6416 ( .B(n5402), .A(n5399), .S(n6259), .Y(n5406) );
  MUX2X1 U6417 ( .B(\Mem[14][18] ), .A(\Mem[15][18] ), .S(n6407), .Y(n5410) );
  MUX2X1 U6418 ( .B(\Mem[12][18] ), .A(\Mem[13][18] ), .S(n6407), .Y(n5409) );
  MUX2X1 U6419 ( .B(\Mem[10][18] ), .A(\Mem[11][18] ), .S(n6407), .Y(n5413) );
  MUX2X1 U6420 ( .B(\Mem[8][18] ), .A(\Mem[9][18] ), .S(n6407), .Y(n5412) );
  MUX2X1 U6421 ( .B(n5411), .A(n5408), .S(n6259), .Y(n5422) );
  MUX2X1 U6422 ( .B(\Mem[6][18] ), .A(\Mem[7][18] ), .S(n6407), .Y(n5416) );
  MUX2X1 U6423 ( .B(\Mem[4][18] ), .A(\Mem[5][18] ), .S(n6407), .Y(n5415) );
  MUX2X1 U6424 ( .B(\Mem[2][18] ), .A(\Mem[3][18] ), .S(n6407), .Y(n5419) );
  MUX2X1 U6425 ( .B(\Mem[0][18] ), .A(\Mem[1][18] ), .S(n6407), .Y(n5418) );
  MUX2X1 U6426 ( .B(n5417), .A(n5414), .S(n6259), .Y(n5421) );
  MUX2X1 U6427 ( .B(n5420), .A(n5405), .S(n6235), .Y(n5423) );
  MUX2X1 U6428 ( .B(\Mem[62][19] ), .A(\Mem[63][19] ), .S(n6408), .Y(n5427) );
  MUX2X1 U6429 ( .B(\Mem[60][19] ), .A(\Mem[61][19] ), .S(n6408), .Y(n5426) );
  MUX2X1 U6430 ( .B(\Mem[58][19] ), .A(\Mem[59][19] ), .S(n6408), .Y(n5430) );
  MUX2X1 U6431 ( .B(\Mem[56][19] ), .A(\Mem[57][19] ), .S(n6408), .Y(n5429) );
  MUX2X1 U6432 ( .B(n5428), .A(n5425), .S(n6260), .Y(n5439) );
  MUX2X1 U6433 ( .B(\Mem[54][19] ), .A(\Mem[55][19] ), .S(n6408), .Y(n5433) );
  MUX2X1 U6434 ( .B(\Mem[52][19] ), .A(\Mem[53][19] ), .S(n6408), .Y(n5432) );
  MUX2X1 U6435 ( .B(\Mem[50][19] ), .A(\Mem[51][19] ), .S(n6408), .Y(n5436) );
  MUX2X1 U6436 ( .B(\Mem[48][19] ), .A(\Mem[49][19] ), .S(n6408), .Y(n5435) );
  MUX2X1 U6437 ( .B(n5434), .A(n5431), .S(n6260), .Y(n5438) );
  MUX2X1 U6438 ( .B(\Mem[46][19] ), .A(\Mem[47][19] ), .S(n6408), .Y(n5442) );
  MUX2X1 U6439 ( .B(\Mem[44][19] ), .A(\Mem[45][19] ), .S(n6408), .Y(n5441) );
  MUX2X1 U6440 ( .B(\Mem[42][19] ), .A(\Mem[43][19] ), .S(n6408), .Y(n5445) );
  MUX2X1 U6441 ( .B(\Mem[40][19] ), .A(\Mem[41][19] ), .S(n6408), .Y(n5444) );
  MUX2X1 U6442 ( .B(n5443), .A(n5440), .S(n6260), .Y(n5454) );
  MUX2X1 U6443 ( .B(\Mem[38][19] ), .A(\Mem[39][19] ), .S(n6408), .Y(n5448) );
  MUX2X1 U6444 ( .B(\Mem[36][19] ), .A(\Mem[37][19] ), .S(n6409), .Y(n5447) );
  MUX2X1 U6445 ( .B(\Mem[34][19] ), .A(\Mem[35][19] ), .S(n6409), .Y(n5451) );
  MUX2X1 U6446 ( .B(\Mem[32][19] ), .A(\Mem[33][19] ), .S(n6409), .Y(n5450) );
  MUX2X1 U6447 ( .B(n5449), .A(n5446), .S(n6260), .Y(n5453) );
  MUX2X1 U6448 ( .B(n5452), .A(n5437), .S(n6236), .Y(n5486) );
  MUX2X1 U6449 ( .B(\Mem[30][19] ), .A(\Mem[31][19] ), .S(n6409), .Y(n5457) );
  MUX2X1 U6450 ( .B(\Mem[28][19] ), .A(\Mem[29][19] ), .S(n6409), .Y(n5456) );
  MUX2X1 U6451 ( .B(\Mem[26][19] ), .A(\Mem[27][19] ), .S(n6409), .Y(n5460) );
  MUX2X1 U6452 ( .B(\Mem[24][19] ), .A(\Mem[25][19] ), .S(n6409), .Y(n5459) );
  MUX2X1 U6453 ( .B(n5458), .A(n5455), .S(n6260), .Y(n5469) );
  MUX2X1 U6454 ( .B(\Mem[22][19] ), .A(\Mem[23][19] ), .S(n6409), .Y(n5463) );
  MUX2X1 U6455 ( .B(\Mem[20][19] ), .A(\Mem[21][19] ), .S(n6409), .Y(n5462) );
  MUX2X1 U6456 ( .B(\Mem[18][19] ), .A(\Mem[19][19] ), .S(n6409), .Y(n5466) );
  MUX2X1 U6457 ( .B(\Mem[16][19] ), .A(\Mem[17][19] ), .S(n6409), .Y(n5465) );
  MUX2X1 U6458 ( .B(n5464), .A(n5461), .S(n6260), .Y(n5468) );
  MUX2X1 U6459 ( .B(\Mem[14][19] ), .A(\Mem[15][19] ), .S(n6409), .Y(n5472) );
  MUX2X1 U6460 ( .B(\Mem[12][19] ), .A(\Mem[13][19] ), .S(n6409), .Y(n5471) );
  MUX2X1 U6461 ( .B(\Mem[10][19] ), .A(\Mem[11][19] ), .S(n6410), .Y(n5475) );
  MUX2X1 U6462 ( .B(\Mem[8][19] ), .A(\Mem[9][19] ), .S(n6410), .Y(n5474) );
  MUX2X1 U6463 ( .B(n5473), .A(n5470), .S(n6260), .Y(n5484) );
  MUX2X1 U6464 ( .B(\Mem[6][19] ), .A(\Mem[7][19] ), .S(n6410), .Y(n5478) );
  MUX2X1 U6465 ( .B(\Mem[4][19] ), .A(\Mem[5][19] ), .S(n6410), .Y(n5477) );
  MUX2X1 U6466 ( .B(\Mem[2][19] ), .A(\Mem[3][19] ), .S(n6410), .Y(n5481) );
  MUX2X1 U6467 ( .B(\Mem[0][19] ), .A(\Mem[1][19] ), .S(n6410), .Y(n5480) );
  MUX2X1 U6468 ( .B(n5479), .A(n5476), .S(n6260), .Y(n5483) );
  MUX2X1 U6469 ( .B(n5482), .A(n5467), .S(n6236), .Y(n5485) );
  MUX2X1 U6470 ( .B(\Mem[62][20] ), .A(\Mem[63][20] ), .S(n6410), .Y(n5489) );
  MUX2X1 U6471 ( .B(\Mem[60][20] ), .A(\Mem[61][20] ), .S(n6410), .Y(n5488) );
  MUX2X1 U6472 ( .B(\Mem[58][20] ), .A(\Mem[59][20] ), .S(n6410), .Y(n5492) );
  MUX2X1 U6473 ( .B(\Mem[56][20] ), .A(\Mem[57][20] ), .S(n6410), .Y(n5491) );
  MUX2X1 U6474 ( .B(n5490), .A(n5487), .S(n6260), .Y(n5501) );
  MUX2X1 U6475 ( .B(\Mem[54][20] ), .A(\Mem[55][20] ), .S(n6410), .Y(n5495) );
  MUX2X1 U6476 ( .B(\Mem[52][20] ), .A(\Mem[53][20] ), .S(n6410), .Y(n5494) );
  MUX2X1 U6477 ( .B(\Mem[50][20] ), .A(\Mem[51][20] ), .S(n6410), .Y(n5498) );
  MUX2X1 U6478 ( .B(\Mem[48][20] ), .A(\Mem[49][20] ), .S(n6411), .Y(n5497) );
  MUX2X1 U6479 ( .B(n5496), .A(n5493), .S(n6260), .Y(n5500) );
  MUX2X1 U6480 ( .B(\Mem[46][20] ), .A(\Mem[47][20] ), .S(n6411), .Y(n5504) );
  MUX2X1 U6481 ( .B(\Mem[44][20] ), .A(\Mem[45][20] ), .S(n6411), .Y(n5503) );
  MUX2X1 U6482 ( .B(\Mem[42][20] ), .A(\Mem[43][20] ), .S(n6411), .Y(n5507) );
  MUX2X1 U6483 ( .B(\Mem[40][20] ), .A(\Mem[41][20] ), .S(n6411), .Y(n5506) );
  MUX2X1 U6484 ( .B(n5505), .A(n5502), .S(n6260), .Y(n5516) );
  MUX2X1 U6485 ( .B(\Mem[38][20] ), .A(\Mem[39][20] ), .S(n6411), .Y(n5510) );
  MUX2X1 U6486 ( .B(\Mem[36][20] ), .A(\Mem[37][20] ), .S(n6411), .Y(n5509) );
  MUX2X1 U6487 ( .B(\Mem[34][20] ), .A(\Mem[35][20] ), .S(n6411), .Y(n5513) );
  MUX2X1 U6488 ( .B(\Mem[32][20] ), .A(\Mem[33][20] ), .S(n6411), .Y(n5512) );
  MUX2X1 U6489 ( .B(n5511), .A(n5508), .S(n6260), .Y(n5515) );
  MUX2X1 U6490 ( .B(n5514), .A(n5499), .S(n6236), .Y(n5548) );
  MUX2X1 U6491 ( .B(\Mem[30][20] ), .A(\Mem[31][20] ), .S(n6411), .Y(n5519) );
  MUX2X1 U6492 ( .B(\Mem[28][20] ), .A(\Mem[29][20] ), .S(n6411), .Y(n5518) );
  MUX2X1 U6493 ( .B(\Mem[26][20] ), .A(\Mem[27][20] ), .S(n6411), .Y(n5522) );
  MUX2X1 U6494 ( .B(\Mem[24][20] ), .A(\Mem[25][20] ), .S(n6411), .Y(n5521) );
  MUX2X1 U6495 ( .B(n5520), .A(n5517), .S(n6260), .Y(n5531) );
  MUX2X1 U6496 ( .B(\Mem[22][20] ), .A(\Mem[23][20] ), .S(n6412), .Y(n5525) );
  MUX2X1 U6497 ( .B(\Mem[20][20] ), .A(\Mem[21][20] ), .S(n6412), .Y(n5524) );
  MUX2X1 U6498 ( .B(\Mem[18][20] ), .A(\Mem[19][20] ), .S(n6412), .Y(n5528) );
  MUX2X1 U6499 ( .B(\Mem[16][20] ), .A(\Mem[17][20] ), .S(n6412), .Y(n5527) );
  MUX2X1 U6500 ( .B(n5526), .A(n5523), .S(n6261), .Y(n5530) );
  MUX2X1 U6501 ( .B(\Mem[14][20] ), .A(\Mem[15][20] ), .S(n6412), .Y(n5534) );
  MUX2X1 U6502 ( .B(\Mem[12][20] ), .A(\Mem[13][20] ), .S(n6412), .Y(n5533) );
  MUX2X1 U6503 ( .B(\Mem[10][20] ), .A(\Mem[11][20] ), .S(n6412), .Y(n5537) );
  MUX2X1 U6504 ( .B(\Mem[8][20] ), .A(\Mem[9][20] ), .S(n6412), .Y(n5536) );
  MUX2X1 U6505 ( .B(n5535), .A(n5532), .S(n6261), .Y(n5546) );
  MUX2X1 U6506 ( .B(\Mem[6][20] ), .A(\Mem[7][20] ), .S(n6412), .Y(n5540) );
  MUX2X1 U6507 ( .B(\Mem[4][20] ), .A(\Mem[5][20] ), .S(n6412), .Y(n5539) );
  MUX2X1 U6508 ( .B(\Mem[2][20] ), .A(\Mem[3][20] ), .S(n6412), .Y(n5543) );
  MUX2X1 U6509 ( .B(\Mem[0][20] ), .A(\Mem[1][20] ), .S(n6412), .Y(n5542) );
  MUX2X1 U6510 ( .B(n5541), .A(n5538), .S(n6261), .Y(n5545) );
  MUX2X1 U6511 ( .B(n5544), .A(n5529), .S(n6236), .Y(n5547) );
  MUX2X1 U6512 ( .B(\Mem[62][21] ), .A(\Mem[63][21] ), .S(n6412), .Y(n5551) );
  MUX2X1 U6513 ( .B(\Mem[60][21] ), .A(\Mem[61][21] ), .S(n6413), .Y(n5550) );
  MUX2X1 U6514 ( .B(\Mem[58][21] ), .A(\Mem[59][21] ), .S(n6413), .Y(n5554) );
  MUX2X1 U6515 ( .B(\Mem[56][21] ), .A(\Mem[57][21] ), .S(n6413), .Y(n5553) );
  MUX2X1 U6516 ( .B(n5552), .A(n5549), .S(n6261), .Y(n5563) );
  MUX2X1 U6517 ( .B(\Mem[54][21] ), .A(\Mem[55][21] ), .S(n6413), .Y(n5557) );
  MUX2X1 U6518 ( .B(\Mem[52][21] ), .A(\Mem[53][21] ), .S(n6413), .Y(n5556) );
  MUX2X1 U6519 ( .B(\Mem[50][21] ), .A(\Mem[51][21] ), .S(n6413), .Y(n5560) );
  MUX2X1 U6520 ( .B(\Mem[48][21] ), .A(\Mem[49][21] ), .S(n6413), .Y(n5559) );
  MUX2X1 U6521 ( .B(n5558), .A(n5555), .S(n6261), .Y(n5562) );
  MUX2X1 U6522 ( .B(\Mem[46][21] ), .A(\Mem[47][21] ), .S(n6413), .Y(n5566) );
  MUX2X1 U6523 ( .B(\Mem[44][21] ), .A(\Mem[45][21] ), .S(n6413), .Y(n5565) );
  MUX2X1 U6524 ( .B(\Mem[42][21] ), .A(\Mem[43][21] ), .S(n6413), .Y(n5569) );
  MUX2X1 U6525 ( .B(\Mem[40][21] ), .A(\Mem[41][21] ), .S(n6413), .Y(n5568) );
  MUX2X1 U6526 ( .B(n5567), .A(n5564), .S(n6261), .Y(n5578) );
  MUX2X1 U6527 ( .B(\Mem[38][21] ), .A(\Mem[39][21] ), .S(n6413), .Y(n5572) );
  MUX2X1 U6528 ( .B(\Mem[36][21] ), .A(\Mem[37][21] ), .S(n6413), .Y(n5571) );
  MUX2X1 U6529 ( .B(\Mem[34][21] ), .A(\Mem[35][21] ), .S(n6414), .Y(n5575) );
  MUX2X1 U6530 ( .B(\Mem[32][21] ), .A(\Mem[33][21] ), .S(n6414), .Y(n5574) );
  MUX2X1 U6531 ( .B(n5573), .A(n5570), .S(n6261), .Y(n5577) );
  MUX2X1 U6532 ( .B(n5576), .A(n5561), .S(n6236), .Y(n5610) );
  MUX2X1 U6533 ( .B(\Mem[30][21] ), .A(\Mem[31][21] ), .S(n6414), .Y(n5581) );
  MUX2X1 U6534 ( .B(\Mem[28][21] ), .A(\Mem[29][21] ), .S(n6414), .Y(n5580) );
  MUX2X1 U6535 ( .B(\Mem[26][21] ), .A(\Mem[27][21] ), .S(n6414), .Y(n5584) );
  MUX2X1 U6536 ( .B(\Mem[24][21] ), .A(\Mem[25][21] ), .S(n6414), .Y(n5583) );
  MUX2X1 U6537 ( .B(n5582), .A(n5579), .S(n6261), .Y(n5593) );
  MUX2X1 U6538 ( .B(\Mem[22][21] ), .A(\Mem[23][21] ), .S(n6414), .Y(n5587) );
  MUX2X1 U6539 ( .B(\Mem[20][21] ), .A(\Mem[21][21] ), .S(n6414), .Y(n5586) );
  MUX2X1 U6540 ( .B(\Mem[18][21] ), .A(\Mem[19][21] ), .S(n6414), .Y(n5590) );
  MUX2X1 U6541 ( .B(\Mem[16][21] ), .A(\Mem[17][21] ), .S(n6414), .Y(n5589) );
  MUX2X1 U6542 ( .B(n5588), .A(n5585), .S(n6261), .Y(n5592) );
  MUX2X1 U6543 ( .B(\Mem[14][21] ), .A(\Mem[15][21] ), .S(n6414), .Y(n5596) );
  MUX2X1 U6544 ( .B(\Mem[12][21] ), .A(\Mem[13][21] ), .S(n6414), .Y(n5595) );
  MUX2X1 U6545 ( .B(\Mem[10][21] ), .A(\Mem[11][21] ), .S(n6414), .Y(n5599) );
  MUX2X1 U6546 ( .B(\Mem[8][21] ), .A(\Mem[9][21] ), .S(n6415), .Y(n5598) );
  MUX2X1 U6547 ( .B(n5597), .A(n5594), .S(n6261), .Y(n5608) );
  MUX2X1 U6548 ( .B(\Mem[6][21] ), .A(\Mem[7][21] ), .S(n6415), .Y(n5602) );
  MUX2X1 U6549 ( .B(\Mem[4][21] ), .A(\Mem[5][21] ), .S(n6415), .Y(n5601) );
  MUX2X1 U6550 ( .B(\Mem[2][21] ), .A(\Mem[3][21] ), .S(n6415), .Y(n5605) );
  MUX2X1 U6551 ( .B(\Mem[0][21] ), .A(\Mem[1][21] ), .S(n6415), .Y(n5604) );
  MUX2X1 U6552 ( .B(n5603), .A(n5600), .S(n6261), .Y(n5607) );
  MUX2X1 U6553 ( .B(n5606), .A(n5591), .S(n6236), .Y(n5609) );
  MUX2X1 U6554 ( .B(\Mem[62][22] ), .A(\Mem[63][22] ), .S(n6415), .Y(n5613) );
  MUX2X1 U6555 ( .B(\Mem[60][22] ), .A(\Mem[61][22] ), .S(n6415), .Y(n5612) );
  MUX2X1 U6556 ( .B(\Mem[58][22] ), .A(\Mem[59][22] ), .S(n6415), .Y(n5616) );
  MUX2X1 U6557 ( .B(\Mem[56][22] ), .A(\Mem[57][22] ), .S(n6415), .Y(n5615) );
  MUX2X1 U6558 ( .B(n5614), .A(n5611), .S(n6261), .Y(n5625) );
  MUX2X1 U6559 ( .B(\Mem[54][22] ), .A(\Mem[55][22] ), .S(n6415), .Y(n5619) );
  MUX2X1 U6560 ( .B(\Mem[52][22] ), .A(\Mem[53][22] ), .S(n6415), .Y(n5618) );
  MUX2X1 U6561 ( .B(\Mem[50][22] ), .A(\Mem[51][22] ), .S(n6415), .Y(n5622) );
  MUX2X1 U6562 ( .B(\Mem[48][22] ), .A(\Mem[49][22] ), .S(n6415), .Y(n5621) );
  MUX2X1 U6563 ( .B(n5620), .A(n5617), .S(n6261), .Y(n5624) );
  MUX2X1 U6564 ( .B(\Mem[46][22] ), .A(\Mem[47][22] ), .S(n6416), .Y(n5628) );
  MUX2X1 U6565 ( .B(\Mem[44][22] ), .A(\Mem[45][22] ), .S(n6416), .Y(n5627) );
  MUX2X1 U6566 ( .B(\Mem[42][22] ), .A(\Mem[43][22] ), .S(n6416), .Y(n5631) );
  MUX2X1 U6567 ( .B(\Mem[40][22] ), .A(\Mem[41][22] ), .S(n6416), .Y(n5630) );
  MUX2X1 U6568 ( .B(n5629), .A(n5626), .S(n6262), .Y(n5640) );
  MUX2X1 U6569 ( .B(\Mem[38][22] ), .A(\Mem[39][22] ), .S(n6416), .Y(n5634) );
  MUX2X1 U6570 ( .B(\Mem[36][22] ), .A(\Mem[37][22] ), .S(n6416), .Y(n5633) );
  MUX2X1 U6571 ( .B(\Mem[34][22] ), .A(\Mem[35][22] ), .S(n6416), .Y(n5637) );
  MUX2X1 U6572 ( .B(\Mem[32][22] ), .A(\Mem[33][22] ), .S(n6416), .Y(n5636) );
  MUX2X1 U6573 ( .B(n5635), .A(n5632), .S(n6262), .Y(n5639) );
  MUX2X1 U6574 ( .B(n5638), .A(n5623), .S(n6236), .Y(n5672) );
  MUX2X1 U6575 ( .B(\Mem[30][22] ), .A(\Mem[31][22] ), .S(n6416), .Y(n5643) );
  MUX2X1 U6576 ( .B(\Mem[28][22] ), .A(\Mem[29][22] ), .S(n6416), .Y(n5642) );
  MUX2X1 U6577 ( .B(\Mem[26][22] ), .A(\Mem[27][22] ), .S(n6416), .Y(n5646) );
  MUX2X1 U6578 ( .B(\Mem[24][22] ), .A(\Mem[25][22] ), .S(n6416), .Y(n5645) );
  MUX2X1 U6579 ( .B(n5644), .A(n5641), .S(n6262), .Y(n5655) );
  MUX2X1 U6580 ( .B(\Mem[22][22] ), .A(\Mem[23][22] ), .S(n6416), .Y(n5649) );
  MUX2X1 U6581 ( .B(\Mem[20][22] ), .A(\Mem[21][22] ), .S(n6417), .Y(n5648) );
  MUX2X1 U6582 ( .B(\Mem[18][22] ), .A(\Mem[19][22] ), .S(n6417), .Y(n5652) );
  MUX2X1 U6583 ( .B(\Mem[16][22] ), .A(\Mem[17][22] ), .S(n6417), .Y(n5651) );
  MUX2X1 U6584 ( .B(n5650), .A(n5647), .S(n6262), .Y(n5654) );
  MUX2X1 U6585 ( .B(\Mem[14][22] ), .A(\Mem[15][22] ), .S(n6417), .Y(n5658) );
  MUX2X1 U6586 ( .B(\Mem[12][22] ), .A(\Mem[13][22] ), .S(n6417), .Y(n5657) );
  MUX2X1 U6587 ( .B(\Mem[10][22] ), .A(\Mem[11][22] ), .S(n6417), .Y(n5661) );
  MUX2X1 U6588 ( .B(\Mem[8][22] ), .A(\Mem[9][22] ), .S(n6417), .Y(n5660) );
  MUX2X1 U6589 ( .B(n5659), .A(n5656), .S(n6262), .Y(n5670) );
  MUX2X1 U6590 ( .B(\Mem[6][22] ), .A(\Mem[7][22] ), .S(n6417), .Y(n5664) );
  MUX2X1 U6591 ( .B(\Mem[4][22] ), .A(\Mem[5][22] ), .S(n6417), .Y(n5663) );
  MUX2X1 U6592 ( .B(\Mem[2][22] ), .A(\Mem[3][22] ), .S(n6417), .Y(n5667) );
  MUX2X1 U6593 ( .B(\Mem[0][22] ), .A(\Mem[1][22] ), .S(n6417), .Y(n5666) );
  MUX2X1 U6594 ( .B(n5665), .A(n5662), .S(n6262), .Y(n5669) );
  MUX2X1 U6595 ( .B(n5668), .A(n5653), .S(n6236), .Y(n5671) );
  MUX2X1 U6596 ( .B(\Mem[62][23] ), .A(\Mem[63][23] ), .S(n6417), .Y(n5675) );
  MUX2X1 U6597 ( .B(\Mem[60][23] ), .A(\Mem[61][23] ), .S(n6417), .Y(n5674) );
  MUX2X1 U6598 ( .B(\Mem[58][23] ), .A(\Mem[59][23] ), .S(n6418), .Y(n5678) );
  MUX2X1 U6599 ( .B(\Mem[56][23] ), .A(\Mem[57][23] ), .S(n6418), .Y(n5677) );
  MUX2X1 U6600 ( .B(n5676), .A(n5673), .S(n6262), .Y(n5687) );
  MUX2X1 U6601 ( .B(\Mem[54][23] ), .A(\Mem[55][23] ), .S(n6418), .Y(n5681) );
  MUX2X1 U6602 ( .B(\Mem[52][23] ), .A(\Mem[53][23] ), .S(n6418), .Y(n5680) );
  MUX2X1 U6603 ( .B(\Mem[50][23] ), .A(\Mem[51][23] ), .S(n6418), .Y(n5684) );
  MUX2X1 U6604 ( .B(\Mem[48][23] ), .A(\Mem[49][23] ), .S(n6418), .Y(n5683) );
  MUX2X1 U6605 ( .B(n5682), .A(n5679), .S(n6262), .Y(n5686) );
  MUX2X1 U6606 ( .B(\Mem[46][23] ), .A(\Mem[47][23] ), .S(n6418), .Y(n5690) );
  MUX2X1 U6607 ( .B(\Mem[44][23] ), .A(\Mem[45][23] ), .S(n6418), .Y(n5689) );
  MUX2X1 U6608 ( .B(\Mem[42][23] ), .A(\Mem[43][23] ), .S(n6418), .Y(n5693) );
  MUX2X1 U6609 ( .B(\Mem[40][23] ), .A(\Mem[41][23] ), .S(n6418), .Y(n5692) );
  MUX2X1 U6610 ( .B(n5691), .A(n5688), .S(n6262), .Y(n5702) );
  MUX2X1 U6611 ( .B(\Mem[38][23] ), .A(\Mem[39][23] ), .S(n6418), .Y(n5696) );
  MUX2X1 U6612 ( .B(\Mem[36][23] ), .A(\Mem[37][23] ), .S(n6418), .Y(n5695) );
  MUX2X1 U6613 ( .B(\Mem[34][23] ), .A(\Mem[35][23] ), .S(n6418), .Y(n5699) );
  MUX2X1 U6614 ( .B(\Mem[32][23] ), .A(\Mem[33][23] ), .S(n6419), .Y(n5698) );
  MUX2X1 U6615 ( .B(n5697), .A(n5694), .S(n6262), .Y(n5701) );
  MUX2X1 U6616 ( .B(n5700), .A(n5685), .S(n6236), .Y(n5734) );
  MUX2X1 U6617 ( .B(\Mem[30][23] ), .A(\Mem[31][23] ), .S(n6419), .Y(n5705) );
  MUX2X1 U6618 ( .B(\Mem[28][23] ), .A(\Mem[29][23] ), .S(n6419), .Y(n5704) );
  MUX2X1 U6619 ( .B(\Mem[26][23] ), .A(\Mem[27][23] ), .S(n6419), .Y(n5708) );
  MUX2X1 U6620 ( .B(\Mem[24][23] ), .A(\Mem[25][23] ), .S(n6419), .Y(n5707) );
  MUX2X1 U6621 ( .B(n5706), .A(n5703), .S(n6262), .Y(n5717) );
  MUX2X1 U6622 ( .B(\Mem[22][23] ), .A(\Mem[23][23] ), .S(n6419), .Y(n5711) );
  MUX2X1 U6623 ( .B(\Mem[20][23] ), .A(\Mem[21][23] ), .S(n6419), .Y(n5710) );
  MUX2X1 U6624 ( .B(\Mem[18][23] ), .A(\Mem[19][23] ), .S(n6419), .Y(n5714) );
  MUX2X1 U6625 ( .B(\Mem[16][23] ), .A(\Mem[17][23] ), .S(n6419), .Y(n5713) );
  MUX2X1 U6626 ( .B(n5712), .A(n5709), .S(n6262), .Y(n5716) );
  MUX2X1 U6627 ( .B(\Mem[14][23] ), .A(\Mem[15][23] ), .S(n6419), .Y(n5720) );
  MUX2X1 U6628 ( .B(\Mem[12][23] ), .A(\Mem[13][23] ), .S(n6419), .Y(n5719) );
  MUX2X1 U6629 ( .B(\Mem[10][23] ), .A(\Mem[11][23] ), .S(n6419), .Y(n5723) );
  MUX2X1 U6630 ( .B(\Mem[8][23] ), .A(\Mem[9][23] ), .S(n6419), .Y(n5722) );
  MUX2X1 U6631 ( .B(n5721), .A(n5718), .S(n6262), .Y(n5732) );
  MUX2X1 U6632 ( .B(\Mem[6][23] ), .A(\Mem[7][23] ), .S(n6420), .Y(n5726) );
  MUX2X1 U6633 ( .B(\Mem[4][23] ), .A(\Mem[5][23] ), .S(n6420), .Y(n5725) );
  MUX2X1 U6634 ( .B(\Mem[2][23] ), .A(\Mem[3][23] ), .S(n6420), .Y(n5729) );
  MUX2X1 U6635 ( .B(\Mem[0][23] ), .A(\Mem[1][23] ), .S(n6420), .Y(n5728) );
  MUX2X1 U6636 ( .B(n5727), .A(n5724), .S(n6263), .Y(n5731) );
  MUX2X1 U6637 ( .B(n5730), .A(n5715), .S(n6236), .Y(n5733) );
  MUX2X1 U6638 ( .B(\Mem[62][24] ), .A(\Mem[63][24] ), .S(n6420), .Y(n5737) );
  MUX2X1 U6639 ( .B(\Mem[60][24] ), .A(\Mem[61][24] ), .S(n6420), .Y(n5736) );
  MUX2X1 U6640 ( .B(\Mem[58][24] ), .A(\Mem[59][24] ), .S(n6420), .Y(n5740) );
  MUX2X1 U6641 ( .B(\Mem[56][24] ), .A(\Mem[57][24] ), .S(n6420), .Y(n5739) );
  MUX2X1 U6642 ( .B(n5738), .A(n5735), .S(n6263), .Y(n5749) );
  MUX2X1 U6643 ( .B(\Mem[54][24] ), .A(\Mem[55][24] ), .S(n6420), .Y(n5743) );
  MUX2X1 U6644 ( .B(\Mem[52][24] ), .A(\Mem[53][24] ), .S(n6420), .Y(n5742) );
  MUX2X1 U6645 ( .B(\Mem[50][24] ), .A(\Mem[51][24] ), .S(n6420), .Y(n5746) );
  MUX2X1 U6646 ( .B(\Mem[48][24] ), .A(\Mem[49][24] ), .S(n6420), .Y(n5745) );
  MUX2X1 U6647 ( .B(n5744), .A(n5741), .S(n6263), .Y(n5748) );
  MUX2X1 U6648 ( .B(\Mem[46][24] ), .A(\Mem[47][24] ), .S(n6420), .Y(n5752) );
  MUX2X1 U6649 ( .B(\Mem[44][24] ), .A(\Mem[45][24] ), .S(n6421), .Y(n5751) );
  MUX2X1 U6650 ( .B(\Mem[42][24] ), .A(\Mem[43][24] ), .S(n6421), .Y(n5755) );
  MUX2X1 U6651 ( .B(\Mem[40][24] ), .A(\Mem[41][24] ), .S(n6421), .Y(n5754) );
  MUX2X1 U6652 ( .B(n5753), .A(n5750), .S(n6263), .Y(n5764) );
  MUX2X1 U6653 ( .B(\Mem[38][24] ), .A(\Mem[39][24] ), .S(n6421), .Y(n5758) );
  MUX2X1 U6654 ( .B(\Mem[36][24] ), .A(\Mem[37][24] ), .S(n6421), .Y(n5757) );
  MUX2X1 U6655 ( .B(\Mem[34][24] ), .A(\Mem[35][24] ), .S(n6421), .Y(n5761) );
  MUX2X1 U6656 ( .B(\Mem[32][24] ), .A(\Mem[33][24] ), .S(n6421), .Y(n5760) );
  MUX2X1 U6657 ( .B(n5759), .A(n5756), .S(n6263), .Y(n5763) );
  MUX2X1 U6658 ( .B(n5762), .A(n5747), .S(n6236), .Y(n5796) );
  MUX2X1 U6659 ( .B(\Mem[30][24] ), .A(\Mem[31][24] ), .S(n6421), .Y(n5767) );
  MUX2X1 U6660 ( .B(\Mem[28][24] ), .A(\Mem[29][24] ), .S(n6421), .Y(n5766) );
  MUX2X1 U6661 ( .B(\Mem[26][24] ), .A(\Mem[27][24] ), .S(n6421), .Y(n5770) );
  MUX2X1 U6662 ( .B(\Mem[24][24] ), .A(\Mem[25][24] ), .S(n6421), .Y(n5769) );
  MUX2X1 U6663 ( .B(n5768), .A(n5765), .S(n6263), .Y(n5779) );
  MUX2X1 U6664 ( .B(\Mem[22][24] ), .A(\Mem[23][24] ), .S(n6421), .Y(n5773) );
  MUX2X1 U6665 ( .B(\Mem[20][24] ), .A(\Mem[21][24] ), .S(n6421), .Y(n5772) );
  MUX2X1 U6666 ( .B(\Mem[18][24] ), .A(\Mem[19][24] ), .S(n6422), .Y(n5776) );
  MUX2X1 U6667 ( .B(\Mem[16][24] ), .A(\Mem[17][24] ), .S(n6422), .Y(n5775) );
  MUX2X1 U6668 ( .B(n5774), .A(n5771), .S(n6263), .Y(n5778) );
  MUX2X1 U6669 ( .B(\Mem[14][24] ), .A(\Mem[15][24] ), .S(n6422), .Y(n5782) );
  MUX2X1 U6670 ( .B(\Mem[12][24] ), .A(\Mem[13][24] ), .S(n6422), .Y(n5781) );
  MUX2X1 U6671 ( .B(\Mem[10][24] ), .A(\Mem[11][24] ), .S(n6422), .Y(n5785) );
  MUX2X1 U6672 ( .B(\Mem[8][24] ), .A(\Mem[9][24] ), .S(n6422), .Y(n5784) );
  MUX2X1 U6673 ( .B(n5783), .A(n5780), .S(n6263), .Y(n5794) );
  MUX2X1 U6674 ( .B(\Mem[6][24] ), .A(\Mem[7][24] ), .S(n6422), .Y(n5788) );
  MUX2X1 U6675 ( .B(\Mem[4][24] ), .A(\Mem[5][24] ), .S(n6422), .Y(n5787) );
  MUX2X1 U6676 ( .B(\Mem[2][24] ), .A(\Mem[3][24] ), .S(n6422), .Y(n5791) );
  MUX2X1 U6677 ( .B(\Mem[0][24] ), .A(\Mem[1][24] ), .S(n6422), .Y(n5790) );
  MUX2X1 U6678 ( .B(n5789), .A(n5786), .S(n6263), .Y(n5793) );
  MUX2X1 U6679 ( .B(n5792), .A(n5777), .S(n6236), .Y(n5795) );
  MUX2X1 U6680 ( .B(\Mem[62][25] ), .A(\Mem[63][25] ), .S(n6422), .Y(n5799) );
  MUX2X1 U6681 ( .B(\Mem[60][25] ), .A(\Mem[61][25] ), .S(n6422), .Y(n5798) );
  MUX2X1 U6682 ( .B(\Mem[58][25] ), .A(\Mem[59][25] ), .S(n6422), .Y(n5802) );
  MUX2X1 U6683 ( .B(\Mem[56][25] ), .A(\Mem[57][25] ), .S(n6423), .Y(n5801) );
  MUX2X1 U6684 ( .B(n5800), .A(n5797), .S(n6263), .Y(n5811) );
  MUX2X1 U6685 ( .B(\Mem[54][25] ), .A(\Mem[55][25] ), .S(n6423), .Y(n5805) );
  MUX2X1 U6686 ( .B(\Mem[52][25] ), .A(\Mem[53][25] ), .S(n6423), .Y(n5804) );
  MUX2X1 U6687 ( .B(\Mem[50][25] ), .A(\Mem[51][25] ), .S(n6423), .Y(n5808) );
  MUX2X1 U6688 ( .B(\Mem[48][25] ), .A(\Mem[49][25] ), .S(n6423), .Y(n5807) );
  MUX2X1 U6689 ( .B(n5806), .A(n5803), .S(n6263), .Y(n5810) );
  MUX2X1 U6690 ( .B(\Mem[46][25] ), .A(\Mem[47][25] ), .S(n6423), .Y(n5814) );
  MUX2X1 U6691 ( .B(\Mem[44][25] ), .A(\Mem[45][25] ), .S(n6423), .Y(n5813) );
  MUX2X1 U6692 ( .B(\Mem[42][25] ), .A(\Mem[43][25] ), .S(n6423), .Y(n5817) );
  MUX2X1 U6693 ( .B(\Mem[40][25] ), .A(\Mem[41][25] ), .S(n6423), .Y(n5816) );
  MUX2X1 U6694 ( .B(n5815), .A(n5812), .S(n6263), .Y(n5826) );
  MUX2X1 U6695 ( .B(\Mem[38][25] ), .A(\Mem[39][25] ), .S(n6423), .Y(n5820) );
  MUX2X1 U6696 ( .B(\Mem[36][25] ), .A(\Mem[37][25] ), .S(n6423), .Y(n5819) );
  MUX2X1 U6697 ( .B(\Mem[34][25] ), .A(\Mem[35][25] ), .S(n6423), .Y(n5823) );
  MUX2X1 U6698 ( .B(\Mem[32][25] ), .A(\Mem[33][25] ), .S(n6423), .Y(n5822) );
  MUX2X1 U6699 ( .B(n5821), .A(n5818), .S(n6263), .Y(n5825) );
  MUX2X1 U6700 ( .B(n5824), .A(n5809), .S(n6236), .Y(n5858) );
  MUX2X1 U6701 ( .B(\Mem[30][25] ), .A(\Mem[31][25] ), .S(n6424), .Y(n5829) );
  MUX2X1 U6702 ( .B(\Mem[28][25] ), .A(\Mem[29][25] ), .S(n6424), .Y(n5828) );
  MUX2X1 U6703 ( .B(\Mem[26][25] ), .A(\Mem[27][25] ), .S(n6424), .Y(n5832) );
  MUX2X1 U6704 ( .B(\Mem[24][25] ), .A(\Mem[25][25] ), .S(n6424), .Y(n5831) );
  MUX2X1 U6705 ( .B(n5830), .A(n5827), .S(n6264), .Y(n5841) );
  MUX2X1 U6706 ( .B(\Mem[22][25] ), .A(\Mem[23][25] ), .S(n6424), .Y(n5835) );
  MUX2X1 U6707 ( .B(\Mem[20][25] ), .A(\Mem[21][25] ), .S(n6424), .Y(n5834) );
  MUX2X1 U6708 ( .B(\Mem[18][25] ), .A(\Mem[19][25] ), .S(n6424), .Y(n5838) );
  MUX2X1 U6709 ( .B(\Mem[16][25] ), .A(\Mem[17][25] ), .S(n6424), .Y(n5837) );
  MUX2X1 U6710 ( .B(n5836), .A(n5833), .S(n6264), .Y(n5840) );
  MUX2X1 U6711 ( .B(\Mem[14][25] ), .A(\Mem[15][25] ), .S(n6424), .Y(n5844) );
  MUX2X1 U6712 ( .B(\Mem[12][25] ), .A(\Mem[13][25] ), .S(n6424), .Y(n5843) );
  MUX2X1 U6713 ( .B(\Mem[10][25] ), .A(\Mem[11][25] ), .S(n6424), .Y(n5847) );
  MUX2X1 U6714 ( .B(\Mem[8][25] ), .A(\Mem[9][25] ), .S(n6424), .Y(n5846) );
  MUX2X1 U6715 ( .B(n5845), .A(n5842), .S(n6264), .Y(n5856) );
  MUX2X1 U6716 ( .B(\Mem[6][25] ), .A(\Mem[7][25] ), .S(n6424), .Y(n5850) );
  MUX2X1 U6717 ( .B(\Mem[4][25] ), .A(\Mem[5][25] ), .S(n6425), .Y(n5849) );
  MUX2X1 U6718 ( .B(\Mem[2][25] ), .A(\Mem[3][25] ), .S(n6425), .Y(n5853) );
  MUX2X1 U6719 ( .B(\Mem[0][25] ), .A(\Mem[1][25] ), .S(n6425), .Y(n5852) );
  MUX2X1 U6720 ( .B(n5851), .A(n5848), .S(n6264), .Y(n5855) );
  MUX2X1 U6721 ( .B(n5854), .A(n5839), .S(n6237), .Y(n5857) );
  MUX2X1 U6722 ( .B(\Mem[62][26] ), .A(\Mem[63][26] ), .S(n6425), .Y(n5861) );
  MUX2X1 U6723 ( .B(\Mem[60][26] ), .A(\Mem[61][26] ), .S(n6425), .Y(n5860) );
  MUX2X1 U6724 ( .B(\Mem[58][26] ), .A(\Mem[59][26] ), .S(n6425), .Y(n5864) );
  MUX2X1 U6725 ( .B(\Mem[56][26] ), .A(\Mem[57][26] ), .S(n6425), .Y(n5863) );
  MUX2X1 U6726 ( .B(n5862), .A(n5859), .S(n6264), .Y(n5873) );
  MUX2X1 U6727 ( .B(\Mem[54][26] ), .A(\Mem[55][26] ), .S(n6425), .Y(n5867) );
  MUX2X1 U6728 ( .B(\Mem[52][26] ), .A(\Mem[53][26] ), .S(n6425), .Y(n5866) );
  MUX2X1 U6729 ( .B(\Mem[50][26] ), .A(\Mem[51][26] ), .S(n6425), .Y(n5870) );
  MUX2X1 U6730 ( .B(\Mem[48][26] ), .A(\Mem[49][26] ), .S(n6425), .Y(n5869) );
  MUX2X1 U6731 ( .B(n5868), .A(n5865), .S(n6264), .Y(n5872) );
  MUX2X1 U6732 ( .B(\Mem[46][26] ), .A(\Mem[47][26] ), .S(n6425), .Y(n5876) );
  MUX2X1 U6733 ( .B(\Mem[44][26] ), .A(\Mem[45][26] ), .S(n6425), .Y(n5875) );
  MUX2X1 U6734 ( .B(\Mem[42][26] ), .A(\Mem[43][26] ), .S(n6426), .Y(n5879) );
  MUX2X1 U6735 ( .B(\Mem[40][26] ), .A(\Mem[41][26] ), .S(n6426), .Y(n5878) );
  MUX2X1 U6736 ( .B(n5877), .A(n5874), .S(n6264), .Y(n5888) );
  MUX2X1 U6737 ( .B(\Mem[38][26] ), .A(\Mem[39][26] ), .S(n6426), .Y(n5882) );
  MUX2X1 U6738 ( .B(\Mem[36][26] ), .A(\Mem[37][26] ), .S(n6426), .Y(n5881) );
  MUX2X1 U6739 ( .B(\Mem[34][26] ), .A(\Mem[35][26] ), .S(n6426), .Y(n5885) );
  MUX2X1 U6740 ( .B(\Mem[32][26] ), .A(\Mem[33][26] ), .S(n6426), .Y(n5884) );
  MUX2X1 U6741 ( .B(n5883), .A(n5880), .S(n6264), .Y(n5887) );
  MUX2X1 U6742 ( .B(n5886), .A(n5871), .S(n6237), .Y(n5920) );
  MUX2X1 U6743 ( .B(\Mem[30][26] ), .A(\Mem[31][26] ), .S(n6426), .Y(n5891) );
  MUX2X1 U6744 ( .B(\Mem[28][26] ), .A(\Mem[29][26] ), .S(n6426), .Y(n5890) );
  MUX2X1 U6745 ( .B(\Mem[26][26] ), .A(\Mem[27][26] ), .S(n6426), .Y(n5894) );
  MUX2X1 U6746 ( .B(\Mem[24][26] ), .A(\Mem[25][26] ), .S(n6426), .Y(n5893) );
  MUX2X1 U6747 ( .B(n5892), .A(n5889), .S(n6264), .Y(n5903) );
  MUX2X1 U6748 ( .B(\Mem[22][26] ), .A(\Mem[23][26] ), .S(n6426), .Y(n5897) );
  MUX2X1 U6749 ( .B(\Mem[20][26] ), .A(\Mem[21][26] ), .S(n6426), .Y(n5896) );
  MUX2X1 U6750 ( .B(\Mem[18][26] ), .A(\Mem[19][26] ), .S(n6426), .Y(n5900) );
  MUX2X1 U6751 ( .B(\Mem[16][26] ), .A(\Mem[17][26] ), .S(n6427), .Y(n5899) );
  MUX2X1 U6752 ( .B(n5898), .A(n5895), .S(n6264), .Y(n5902) );
  MUX2X1 U6753 ( .B(\Mem[14][26] ), .A(\Mem[15][26] ), .S(n6427), .Y(n5906) );
  MUX2X1 U6754 ( .B(\Mem[12][26] ), .A(\Mem[13][26] ), .S(n6427), .Y(n5905) );
  MUX2X1 U6755 ( .B(\Mem[10][26] ), .A(\Mem[11][26] ), .S(n6427), .Y(n5909) );
  MUX2X1 U6756 ( .B(\Mem[8][26] ), .A(\Mem[9][26] ), .S(n6427), .Y(n5908) );
  MUX2X1 U6757 ( .B(n5907), .A(n5904), .S(n6264), .Y(n5918) );
  MUX2X1 U6758 ( .B(\Mem[6][26] ), .A(\Mem[7][26] ), .S(n6427), .Y(n5912) );
  MUX2X1 U6759 ( .B(\Mem[4][26] ), .A(\Mem[5][26] ), .S(n6427), .Y(n5911) );
  MUX2X1 U6760 ( .B(\Mem[2][26] ), .A(\Mem[3][26] ), .S(n6427), .Y(n5915) );
  MUX2X1 U6761 ( .B(\Mem[0][26] ), .A(\Mem[1][26] ), .S(n6427), .Y(n5914) );
  MUX2X1 U6762 ( .B(n5913), .A(n5910), .S(n6264), .Y(n5917) );
  MUX2X1 U6763 ( .B(n5916), .A(n5901), .S(n6237), .Y(n5919) );
  MUX2X1 U6764 ( .B(\Mem[62][27] ), .A(\Mem[63][27] ), .S(n6427), .Y(n5923) );
  MUX2X1 U6765 ( .B(\Mem[60][27] ), .A(\Mem[61][27] ), .S(n6427), .Y(n5922) );
  MUX2X1 U6766 ( .B(\Mem[58][27] ), .A(\Mem[59][27] ), .S(n6427), .Y(n5926) );
  MUX2X1 U6767 ( .B(\Mem[56][27] ), .A(\Mem[57][27] ), .S(n6427), .Y(n5925) );
  MUX2X1 U6768 ( .B(n5924), .A(n5921), .S(n6264), .Y(n5935) );
  MUX2X1 U6769 ( .B(\Mem[54][27] ), .A(\Mem[55][27] ), .S(n6428), .Y(n5929) );
  MUX2X1 U6770 ( .B(\Mem[52][27] ), .A(\Mem[53][27] ), .S(n6428), .Y(n5928) );
  MUX2X1 U6771 ( .B(\Mem[50][27] ), .A(\Mem[51][27] ), .S(n6428), .Y(n5932) );
  MUX2X1 U6772 ( .B(\Mem[48][27] ), .A(\Mem[49][27] ), .S(n6428), .Y(n5931) );
  MUX2X1 U6773 ( .B(n5930), .A(n5927), .S(n6265), .Y(n5934) );
  MUX2X1 U6774 ( .B(\Mem[46][27] ), .A(\Mem[47][27] ), .S(n6428), .Y(n5938) );
  MUX2X1 U6775 ( .B(\Mem[44][27] ), .A(\Mem[45][27] ), .S(n6428), .Y(n5937) );
  MUX2X1 U6776 ( .B(\Mem[42][27] ), .A(\Mem[43][27] ), .S(n6428), .Y(n5941) );
  MUX2X1 U6777 ( .B(\Mem[40][27] ), .A(\Mem[41][27] ), .S(n6428), .Y(n5940) );
  MUX2X1 U6778 ( .B(n5939), .A(n5936), .S(n6265), .Y(n5950) );
  MUX2X1 U6779 ( .B(\Mem[38][27] ), .A(\Mem[39][27] ), .S(n6428), .Y(n5944) );
  MUX2X1 U6780 ( .B(\Mem[36][27] ), .A(\Mem[37][27] ), .S(n6428), .Y(n5943) );
  MUX2X1 U6781 ( .B(\Mem[34][27] ), .A(\Mem[35][27] ), .S(n6428), .Y(n5947) );
  MUX2X1 U6782 ( .B(\Mem[32][27] ), .A(\Mem[33][27] ), .S(n6428), .Y(n5946) );
  MUX2X1 U6783 ( .B(n5945), .A(n5942), .S(n6265), .Y(n5949) );
  MUX2X1 U6784 ( .B(n5948), .A(n5933), .S(n6237), .Y(n5982) );
  MUX2X1 U6785 ( .B(\Mem[30][27] ), .A(\Mem[31][27] ), .S(n6428), .Y(n5953) );
  MUX2X1 U6786 ( .B(\Mem[28][27] ), .A(\Mem[29][27] ), .S(n6429), .Y(n5952) );
  MUX2X1 U6787 ( .B(\Mem[26][27] ), .A(\Mem[27][27] ), .S(n6429), .Y(n5956) );
  MUX2X1 U6788 ( .B(\Mem[24][27] ), .A(\Mem[25][27] ), .S(n6429), .Y(n5955) );
  MUX2X1 U6789 ( .B(n5954), .A(n5951), .S(n6265), .Y(n5965) );
  MUX2X1 U6790 ( .B(\Mem[22][27] ), .A(\Mem[23][27] ), .S(n6429), .Y(n5959) );
  MUX2X1 U6791 ( .B(\Mem[20][27] ), .A(\Mem[21][27] ), .S(n6429), .Y(n5958) );
  MUX2X1 U6792 ( .B(\Mem[18][27] ), .A(\Mem[19][27] ), .S(n6429), .Y(n5962) );
  MUX2X1 U6793 ( .B(\Mem[16][27] ), .A(\Mem[17][27] ), .S(n6429), .Y(n5961) );
  MUX2X1 U6794 ( .B(n5960), .A(n5957), .S(n6265), .Y(n5964) );
  MUX2X1 U6795 ( .B(\Mem[14][27] ), .A(\Mem[15][27] ), .S(n6429), .Y(n5968) );
  MUX2X1 U6796 ( .B(\Mem[12][27] ), .A(\Mem[13][27] ), .S(n6429), .Y(n5967) );
  MUX2X1 U6797 ( .B(\Mem[10][27] ), .A(\Mem[11][27] ), .S(n6429), .Y(n5971) );
  MUX2X1 U6798 ( .B(\Mem[8][27] ), .A(\Mem[9][27] ), .S(n6429), .Y(n5970) );
  MUX2X1 U6799 ( .B(n5969), .A(n5966), .S(n6265), .Y(n5980) );
  MUX2X1 U6800 ( .B(\Mem[6][27] ), .A(\Mem[7][27] ), .S(n6429), .Y(n5974) );
  MUX2X1 U6801 ( .B(\Mem[4][27] ), .A(\Mem[5][27] ), .S(n6429), .Y(n5973) );
  MUX2X1 U6802 ( .B(\Mem[2][27] ), .A(\Mem[3][27] ), .S(n6430), .Y(n5977) );
  MUX2X1 U6803 ( .B(\Mem[0][27] ), .A(\Mem[1][27] ), .S(n6430), .Y(n5976) );
  MUX2X1 U6804 ( .B(n5975), .A(n5972), .S(n6265), .Y(n5979) );
  MUX2X1 U6805 ( .B(n5978), .A(n5963), .S(n6237), .Y(n5981) );
  MUX2X1 U6806 ( .B(\Mem[62][28] ), .A(\Mem[63][28] ), .S(n6430), .Y(n5985) );
  MUX2X1 U6807 ( .B(\Mem[60][28] ), .A(\Mem[61][28] ), .S(n6430), .Y(n5984) );
  MUX2X1 U6808 ( .B(\Mem[58][28] ), .A(\Mem[59][28] ), .S(n6430), .Y(n5988) );
  MUX2X1 U6809 ( .B(\Mem[56][28] ), .A(\Mem[57][28] ), .S(n6430), .Y(n5987) );
  MUX2X1 U6810 ( .B(n5986), .A(n5983), .S(n6265), .Y(n5997) );
  MUX2X1 U6811 ( .B(\Mem[54][28] ), .A(\Mem[55][28] ), .S(n6430), .Y(n5991) );
  MUX2X1 U6812 ( .B(\Mem[52][28] ), .A(\Mem[53][28] ), .S(n6430), .Y(n5990) );
  MUX2X1 U6813 ( .B(\Mem[50][28] ), .A(\Mem[51][28] ), .S(n6430), .Y(n5994) );
  MUX2X1 U6814 ( .B(\Mem[48][28] ), .A(\Mem[49][28] ), .S(n6430), .Y(n5993) );
  MUX2X1 U6815 ( .B(n5992), .A(n5989), .S(n6265), .Y(n5996) );
  MUX2X1 U6816 ( .B(\Mem[46][28] ), .A(\Mem[47][28] ), .S(n6430), .Y(n6000) );
  MUX2X1 U6817 ( .B(\Mem[44][28] ), .A(\Mem[45][28] ), .S(n6430), .Y(n5999) );
  MUX2X1 U6818 ( .B(\Mem[42][28] ), .A(\Mem[43][28] ), .S(n6430), .Y(n6003) );
  MUX2X1 U6819 ( .B(\Mem[40][28] ), .A(\Mem[41][28] ), .S(n6431), .Y(n6002) );
  MUX2X1 U6820 ( .B(n6001), .A(n5998), .S(n6265), .Y(n6012) );
  MUX2X1 U6821 ( .B(\Mem[38][28] ), .A(\Mem[39][28] ), .S(n6431), .Y(n6006) );
  MUX2X1 U6822 ( .B(\Mem[36][28] ), .A(\Mem[37][28] ), .S(n6431), .Y(n6005) );
  MUX2X1 U6823 ( .B(\Mem[34][28] ), .A(\Mem[35][28] ), .S(n6431), .Y(n6009) );
  MUX2X1 U6824 ( .B(\Mem[32][28] ), .A(\Mem[33][28] ), .S(n6431), .Y(n6008) );
  MUX2X1 U6825 ( .B(n6007), .A(n6004), .S(n6265), .Y(n6011) );
  MUX2X1 U6826 ( .B(n6010), .A(n5995), .S(n6237), .Y(n6044) );
  MUX2X1 U6827 ( .B(\Mem[30][28] ), .A(\Mem[31][28] ), .S(n6431), .Y(n6015) );
  MUX2X1 U6828 ( .B(\Mem[28][28] ), .A(\Mem[29][28] ), .S(n6431), .Y(n6014) );
  MUX2X1 U6829 ( .B(\Mem[26][28] ), .A(\Mem[27][28] ), .S(n6431), .Y(n6018) );
  MUX2X1 U6830 ( .B(\Mem[24][28] ), .A(\Mem[25][28] ), .S(n6431), .Y(n6017) );
  MUX2X1 U6831 ( .B(n6016), .A(n6013), .S(n6265), .Y(n6027) );
  MUX2X1 U6832 ( .B(\Mem[22][28] ), .A(\Mem[23][28] ), .S(n6431), .Y(n6021) );
  MUX2X1 U6833 ( .B(\Mem[20][28] ), .A(\Mem[21][28] ), .S(n6431), .Y(n6020) );
  MUX2X1 U6834 ( .B(\Mem[18][28] ), .A(\Mem[19][28] ), .S(n6431), .Y(n6024) );
  MUX2X1 U6835 ( .B(\Mem[16][28] ), .A(\Mem[17][28] ), .S(n6431), .Y(n6023) );
  MUX2X1 U6836 ( .B(n6022), .A(n6019), .S(n6265), .Y(n6026) );
  MUX2X1 U6837 ( .B(\Mem[14][28] ), .A(\Mem[15][28] ), .S(n6432), .Y(n6030) );
  MUX2X1 U6838 ( .B(\Mem[12][28] ), .A(\Mem[13][28] ), .S(n6432), .Y(n6029) );
  MUX2X1 U6839 ( .B(\Mem[10][28] ), .A(\Mem[11][28] ), .S(n6432), .Y(n6033) );
  MUX2X1 U6840 ( .B(\Mem[8][28] ), .A(\Mem[9][28] ), .S(n6432), .Y(n6032) );
  MUX2X1 U6841 ( .B(n6031), .A(n6028), .S(n6266), .Y(n6042) );
  MUX2X1 U6842 ( .B(\Mem[6][28] ), .A(\Mem[7][28] ), .S(n6432), .Y(n6036) );
  MUX2X1 U6843 ( .B(\Mem[4][28] ), .A(\Mem[5][28] ), .S(n6432), .Y(n6035) );
  MUX2X1 U6844 ( .B(\Mem[2][28] ), .A(\Mem[3][28] ), .S(n6432), .Y(n6039) );
  MUX2X1 U6845 ( .B(\Mem[0][28] ), .A(\Mem[1][28] ), .S(n6432), .Y(n6038) );
  MUX2X1 U6846 ( .B(n6037), .A(n6034), .S(n6266), .Y(n6041) );
  MUX2X1 U6847 ( .B(n6040), .A(n6025), .S(n6237), .Y(n6043) );
  MUX2X1 U6848 ( .B(\Mem[62][29] ), .A(\Mem[63][29] ), .S(n6432), .Y(n6047) );
  MUX2X1 U6849 ( .B(\Mem[60][29] ), .A(\Mem[61][29] ), .S(n6432), .Y(n6046) );
  MUX2X1 U6850 ( .B(\Mem[58][29] ), .A(\Mem[59][29] ), .S(n6432), .Y(n6050) );
  MUX2X1 U6851 ( .B(\Mem[56][29] ), .A(\Mem[57][29] ), .S(n6432), .Y(n6049) );
  MUX2X1 U6852 ( .B(n6048), .A(n6045), .S(n6266), .Y(n6059) );
  MUX2X1 U6853 ( .B(\Mem[54][29] ), .A(\Mem[55][29] ), .S(n6432), .Y(n6053) );
  MUX2X1 U6854 ( .B(\Mem[52][29] ), .A(\Mem[53][29] ), .S(n6433), .Y(n6052) );
  MUX2X1 U6855 ( .B(\Mem[50][29] ), .A(\Mem[51][29] ), .S(n6433), .Y(n6056) );
  MUX2X1 U6856 ( .B(\Mem[48][29] ), .A(\Mem[49][29] ), .S(n6433), .Y(n6055) );
  MUX2X1 U6857 ( .B(n6054), .A(n6051), .S(n6266), .Y(n6058) );
  MUX2X1 U6858 ( .B(\Mem[46][29] ), .A(\Mem[47][29] ), .S(n6433), .Y(n6062) );
  MUX2X1 U6859 ( .B(\Mem[44][29] ), .A(\Mem[45][29] ), .S(n6433), .Y(n6061) );
  MUX2X1 U6860 ( .B(\Mem[42][29] ), .A(\Mem[43][29] ), .S(n6433), .Y(n6065) );
  MUX2X1 U6861 ( .B(\Mem[40][29] ), .A(\Mem[41][29] ), .S(n6433), .Y(n6064) );
  MUX2X1 U6862 ( .B(n6063), .A(n6060), .S(n6266), .Y(n6074) );
  MUX2X1 U6863 ( .B(\Mem[38][29] ), .A(\Mem[39][29] ), .S(n6433), .Y(n6068) );
  MUX2X1 U6864 ( .B(\Mem[36][29] ), .A(\Mem[37][29] ), .S(n6433), .Y(n6067) );
  MUX2X1 U6865 ( .B(\Mem[34][29] ), .A(\Mem[35][29] ), .S(n6433), .Y(n6071) );
  MUX2X1 U6866 ( .B(\Mem[32][29] ), .A(\Mem[33][29] ), .S(n6433), .Y(n6070) );
  MUX2X1 U6867 ( .B(n6069), .A(n6066), .S(n6266), .Y(n6073) );
  MUX2X1 U6868 ( .B(n6072), .A(n6057), .S(n6237), .Y(n6106) );
  MUX2X1 U6869 ( .B(\Mem[30][29] ), .A(\Mem[31][29] ), .S(n6433), .Y(n6077) );
  MUX2X1 U6870 ( .B(\Mem[28][29] ), .A(\Mem[29][29] ), .S(n6433), .Y(n6076) );
  MUX2X1 U6871 ( .B(\Mem[26][29] ), .A(\Mem[27][29] ), .S(n6434), .Y(n6080) );
  MUX2X1 U6872 ( .B(\Mem[24][29] ), .A(\Mem[25][29] ), .S(n6434), .Y(n6079) );
  MUX2X1 U6873 ( .B(n6078), .A(n6075), .S(n6266), .Y(n6089) );
  MUX2X1 U6874 ( .B(\Mem[22][29] ), .A(\Mem[23][29] ), .S(n6434), .Y(n6083) );
  MUX2X1 U6875 ( .B(\Mem[20][29] ), .A(\Mem[21][29] ), .S(n6434), .Y(n6082) );
  MUX2X1 U6876 ( .B(\Mem[18][29] ), .A(\Mem[19][29] ), .S(n6434), .Y(n6086) );
  MUX2X1 U6877 ( .B(\Mem[16][29] ), .A(\Mem[17][29] ), .S(n6434), .Y(n6085) );
  MUX2X1 U6878 ( .B(n6084), .A(n6081), .S(n6266), .Y(n6088) );
  MUX2X1 U6879 ( .B(\Mem[14][29] ), .A(\Mem[15][29] ), .S(n6434), .Y(n6092) );
  MUX2X1 U6880 ( .B(\Mem[12][29] ), .A(\Mem[13][29] ), .S(n6434), .Y(n6091) );
  MUX2X1 U6881 ( .B(\Mem[10][29] ), .A(\Mem[11][29] ), .S(n6434), .Y(n6095) );
  MUX2X1 U6882 ( .B(\Mem[8][29] ), .A(\Mem[9][29] ), .S(n6434), .Y(n6094) );
  MUX2X1 U6883 ( .B(n6093), .A(n6090), .S(n6266), .Y(n6104) );
  MUX2X1 U6884 ( .B(\Mem[6][29] ), .A(\Mem[7][29] ), .S(n6434), .Y(n6098) );
  MUX2X1 U6885 ( .B(\Mem[4][29] ), .A(\Mem[5][29] ), .S(n6434), .Y(n6097) );
  MUX2X1 U6886 ( .B(\Mem[2][29] ), .A(\Mem[3][29] ), .S(n6434), .Y(n6101) );
  MUX2X1 U6887 ( .B(\Mem[0][29] ), .A(\Mem[1][29] ), .S(n6435), .Y(n6100) );
  MUX2X1 U6888 ( .B(n6099), .A(n6096), .S(n6266), .Y(n6103) );
  MUX2X1 U6889 ( .B(n6102), .A(n6087), .S(n6237), .Y(n6105) );
  MUX2X1 U6890 ( .B(\Mem[62][30] ), .A(\Mem[63][30] ), .S(n6435), .Y(n6109) );
  MUX2X1 U6891 ( .B(\Mem[60][30] ), .A(\Mem[61][30] ), .S(n6435), .Y(n6108) );
  MUX2X1 U6892 ( .B(\Mem[58][30] ), .A(\Mem[59][30] ), .S(n6435), .Y(n6112) );
  MUX2X1 U6893 ( .B(\Mem[56][30] ), .A(\Mem[57][30] ), .S(n6435), .Y(n6111) );
  MUX2X1 U6894 ( .B(n6110), .A(n6107), .S(n6266), .Y(n6121) );
  MUX2X1 U6895 ( .B(\Mem[54][30] ), .A(\Mem[55][30] ), .S(n6435), .Y(n6115) );
  MUX2X1 U6896 ( .B(\Mem[52][30] ), .A(\Mem[53][30] ), .S(n6435), .Y(n6114) );
  MUX2X1 U6897 ( .B(\Mem[50][30] ), .A(\Mem[51][30] ), .S(n6435), .Y(n6118) );
  MUX2X1 U6898 ( .B(\Mem[48][30] ), .A(\Mem[49][30] ), .S(n6435), .Y(n6117) );
  MUX2X1 U6899 ( .B(n6116), .A(n6113), .S(n6266), .Y(n6120) );
  MUX2X1 U6900 ( .B(\Mem[46][30] ), .A(\Mem[47][30] ), .S(n6435), .Y(n6124) );
  MUX2X1 U6901 ( .B(\Mem[44][30] ), .A(\Mem[45][30] ), .S(n6435), .Y(n6123) );
  MUX2X1 U6902 ( .B(\Mem[42][30] ), .A(\Mem[43][30] ), .S(n6435), .Y(n6127) );
  MUX2X1 U6903 ( .B(\Mem[40][30] ), .A(\Mem[41][30] ), .S(n6435), .Y(n6126) );
  MUX2X1 U6904 ( .B(n6125), .A(n6122), .S(n6266), .Y(n6136) );
  MUX2X1 U6905 ( .B(\Mem[38][30] ), .A(\Mem[39][30] ), .S(n6436), .Y(n6130) );
  MUX2X1 U6906 ( .B(\Mem[36][30] ), .A(\Mem[37][30] ), .S(n6436), .Y(n6129) );
  MUX2X1 U6907 ( .B(\Mem[34][30] ), .A(\Mem[35][30] ), .S(n6436), .Y(n6133) );
  MUX2X1 U6908 ( .B(\Mem[32][30] ), .A(\Mem[33][30] ), .S(n6436), .Y(n6132) );
  MUX2X1 U6909 ( .B(n6131), .A(n6128), .S(n6267), .Y(n6135) );
  MUX2X1 U6910 ( .B(n6134), .A(n6119), .S(n6237), .Y(n6168) );
  MUX2X1 U6911 ( .B(\Mem[30][30] ), .A(\Mem[31][30] ), .S(n6436), .Y(n6139) );
  MUX2X1 U6912 ( .B(\Mem[28][30] ), .A(\Mem[29][30] ), .S(n6436), .Y(n6138) );
  MUX2X1 U6913 ( .B(\Mem[26][30] ), .A(\Mem[27][30] ), .S(n6436), .Y(n6142) );
  MUX2X1 U6914 ( .B(\Mem[24][30] ), .A(\Mem[25][30] ), .S(n6436), .Y(n6141) );
  MUX2X1 U6915 ( .B(n6140), .A(n6137), .S(n6267), .Y(n6151) );
  MUX2X1 U6916 ( .B(\Mem[22][30] ), .A(\Mem[23][30] ), .S(n6436), .Y(n6145) );
  MUX2X1 U6917 ( .B(\Mem[20][30] ), .A(\Mem[21][30] ), .S(n6436), .Y(n6144) );
  MUX2X1 U6918 ( .B(\Mem[18][30] ), .A(\Mem[19][30] ), .S(n6436), .Y(n6148) );
  MUX2X1 U6919 ( .B(\Mem[16][30] ), .A(\Mem[17][30] ), .S(n6436), .Y(n6147) );
  MUX2X1 U6920 ( .B(n6146), .A(n6143), .S(n6267), .Y(n6150) );
  MUX2X1 U6921 ( .B(\Mem[14][30] ), .A(\Mem[15][30] ), .S(n6436), .Y(n6154) );
  MUX2X1 U6922 ( .B(\Mem[12][30] ), .A(\Mem[13][30] ), .S(n6437), .Y(n6153) );
  MUX2X1 U6923 ( .B(\Mem[10][30] ), .A(\Mem[11][30] ), .S(n6437), .Y(n6157) );
  MUX2X1 U6924 ( .B(\Mem[8][30] ), .A(\Mem[9][30] ), .S(n6437), .Y(n6156) );
  MUX2X1 U6925 ( .B(n6155), .A(n6152), .S(n6267), .Y(n6166) );
  MUX2X1 U6926 ( .B(\Mem[6][30] ), .A(\Mem[7][30] ), .S(n6437), .Y(n6160) );
  MUX2X1 U6927 ( .B(\Mem[4][30] ), .A(\Mem[5][30] ), .S(n6437), .Y(n6159) );
  MUX2X1 U6928 ( .B(\Mem[2][30] ), .A(\Mem[3][30] ), .S(n6437), .Y(n6163) );
  MUX2X1 U6929 ( .B(\Mem[0][30] ), .A(\Mem[1][30] ), .S(n6437), .Y(n6162) );
  MUX2X1 U6930 ( .B(n6161), .A(n6158), .S(n6267), .Y(n6165) );
  MUX2X1 U6931 ( .B(n6164), .A(n6149), .S(n6237), .Y(n6167) );
  MUX2X1 U6932 ( .B(\Mem[62][31] ), .A(\Mem[63][31] ), .S(n6437), .Y(n6171) );
  MUX2X1 U6933 ( .B(\Mem[60][31] ), .A(\Mem[61][31] ), .S(n6437), .Y(n6170) );
  MUX2X1 U6934 ( .B(\Mem[58][31] ), .A(\Mem[59][31] ), .S(n6437), .Y(n6174) );
  MUX2X1 U6935 ( .B(\Mem[56][31] ), .A(\Mem[57][31] ), .S(n6437), .Y(n6173) );
  MUX2X1 U6936 ( .B(n6172), .A(n6169), .S(n6267), .Y(n6183) );
  MUX2X1 U6937 ( .B(\Mem[54][31] ), .A(\Mem[55][31] ), .S(n6437), .Y(n6177) );
  MUX2X1 U6938 ( .B(\Mem[52][31] ), .A(\Mem[53][31] ), .S(n6437), .Y(n6176) );
  MUX2X1 U6939 ( .B(\Mem[50][31] ), .A(\Mem[51][31] ), .S(n6438), .Y(n6180) );
  MUX2X1 U6940 ( .B(\Mem[48][31] ), .A(\Mem[49][31] ), .S(n6438), .Y(n6179) );
  MUX2X1 U6941 ( .B(n6178), .A(n6175), .S(n6267), .Y(n6182) );
  MUX2X1 U6942 ( .B(\Mem[46][31] ), .A(\Mem[47][31] ), .S(n6438), .Y(n6186) );
  MUX2X1 U6943 ( .B(\Mem[44][31] ), .A(\Mem[45][31] ), .S(n6438), .Y(n6185) );
  MUX2X1 U6944 ( .B(\Mem[42][31] ), .A(\Mem[43][31] ), .S(n6438), .Y(n6189) );
  MUX2X1 U6945 ( .B(\Mem[40][31] ), .A(\Mem[41][31] ), .S(n6438), .Y(n6188) );
  MUX2X1 U6946 ( .B(n6187), .A(n6184), .S(n6267), .Y(n6198) );
  MUX2X1 U6947 ( .B(\Mem[38][31] ), .A(\Mem[39][31] ), .S(n6438), .Y(n6192) );
  MUX2X1 U6948 ( .B(\Mem[36][31] ), .A(\Mem[37][31] ), .S(n6438), .Y(n6191) );
  MUX2X1 U6949 ( .B(\Mem[34][31] ), .A(\Mem[35][31] ), .S(n6438), .Y(n6195) );
  MUX2X1 U6950 ( .B(\Mem[32][31] ), .A(\Mem[33][31] ), .S(n6438), .Y(n6194) );
  MUX2X1 U6951 ( .B(n6193), .A(n6190), .S(n6267), .Y(n6197) );
  MUX2X1 U6952 ( .B(n6196), .A(n6181), .S(n6237), .Y(n6230) );
  MUX2X1 U6953 ( .B(\Mem[30][31] ), .A(\Mem[31][31] ), .S(n6438), .Y(n6201) );
  MUX2X1 U6954 ( .B(\Mem[28][31] ), .A(\Mem[29][31] ), .S(n6438), .Y(n6200) );
  MUX2X1 U6955 ( .B(\Mem[26][31] ), .A(\Mem[27][31] ), .S(n6438), .Y(n6204) );
  MUX2X1 U6956 ( .B(\Mem[24][31] ), .A(\Mem[25][31] ), .S(n6439), .Y(n6203) );
  MUX2X1 U6957 ( .B(n6202), .A(n6199), .S(n6267), .Y(n6213) );
  MUX2X1 U6958 ( .B(\Mem[22][31] ), .A(\Mem[23][31] ), .S(n6439), .Y(n6207) );
  MUX2X1 U6959 ( .B(\Mem[20][31] ), .A(\Mem[21][31] ), .S(n6439), .Y(n6206) );
  MUX2X1 U6960 ( .B(\Mem[18][31] ), .A(\Mem[19][31] ), .S(n6439), .Y(n6210) );
  MUX2X1 U6961 ( .B(\Mem[16][31] ), .A(\Mem[17][31] ), .S(n6439), .Y(n6209) );
  MUX2X1 U6962 ( .B(n6208), .A(n6205), .S(n6267), .Y(n6212) );
  MUX2X1 U6963 ( .B(\Mem[14][31] ), .A(\Mem[15][31] ), .S(n6439), .Y(n6216) );
  MUX2X1 U6964 ( .B(\Mem[12][31] ), .A(\Mem[13][31] ), .S(n6439), .Y(n6215) );
  MUX2X1 U6965 ( .B(\Mem[10][31] ), .A(\Mem[11][31] ), .S(n6439), .Y(n6219) );
  MUX2X1 U6966 ( .B(\Mem[8][31] ), .A(\Mem[9][31] ), .S(n6439), .Y(n6218) );
  MUX2X1 U6967 ( .B(n6217), .A(n6214), .S(n6267), .Y(n6228) );
  MUX2X1 U6968 ( .B(\Mem[6][31] ), .A(\Mem[7][31] ), .S(n6439), .Y(n6222) );
  MUX2X1 U6969 ( .B(\Mem[4][31] ), .A(\Mem[5][31] ), .S(n6439), .Y(n6221) );
  MUX2X1 U6970 ( .B(\Mem[2][31] ), .A(\Mem[3][31] ), .S(n6439), .Y(n6225) );
  MUX2X1 U6971 ( .B(\Mem[0][31] ), .A(\Mem[1][31] ), .S(n6439), .Y(n6224) );
  MUX2X1 U6972 ( .B(n6223), .A(n6220), .S(n6267), .Y(n6227) );
  MUX2X1 U6973 ( .B(n6226), .A(n6211), .S(n6237), .Y(n6229) );
  INVX2 U6974 ( .A(n1990), .Y(n6940) );
  INVX2 U6975 ( .A(n1989), .Y(n6941) );
  INVX2 U6976 ( .A(n1988), .Y(n6942) );
  INVX2 U6977 ( .A(n1987), .Y(n6943) );
  INVX2 U6978 ( .A(n1986), .Y(n6944) );
  INVX2 U6979 ( .A(n1985), .Y(n6945) );
  INVX2 U6980 ( .A(n1984), .Y(n6946) );
  INVX2 U6981 ( .A(n1983), .Y(n6947) );
  INVX2 U6982 ( .A(n1982), .Y(n6948) );
  INVX2 U6983 ( .A(n1981), .Y(n6949) );
  INVX2 U6984 ( .A(n1980), .Y(n6950) );
  INVX2 U6985 ( .A(n1979), .Y(n6951) );
  INVX2 U6986 ( .A(n1978), .Y(n6952) );
  INVX2 U6987 ( .A(n1977), .Y(n6953) );
  INVX2 U6988 ( .A(n1976), .Y(n6954) );
  INVX2 U6989 ( .A(n1975), .Y(n6955) );
  INVX2 U6990 ( .A(n1974), .Y(n6956) );
  INVX2 U6991 ( .A(n1973), .Y(n6957) );
  INVX2 U6992 ( .A(n1972), .Y(n6958) );
  INVX2 U6993 ( .A(n1971), .Y(n6959) );
  INVX2 U6994 ( .A(n1970), .Y(n6960) );
  INVX2 U6995 ( .A(n1969), .Y(n6961) );
  INVX2 U6996 ( .A(n1968), .Y(n6962) );
  INVX2 U6997 ( .A(n1967), .Y(n6963) );
  INVX2 U6998 ( .A(n1966), .Y(n6964) );
  INVX2 U6999 ( .A(n1965), .Y(n6965) );
  INVX2 U7000 ( .A(n1964), .Y(n6966) );
  INVX2 U7001 ( .A(n1963), .Y(n6967) );
  INVX2 U7002 ( .A(n1962), .Y(n6968) );
  INVX2 U7003 ( .A(n1961), .Y(n6969) );
  INVX2 U7004 ( .A(n1960), .Y(n6970) );
  INVX2 U7005 ( .A(n1958), .Y(n6971) );
  INVX2 U7006 ( .A(DIN[9]), .Y(n6972) );
  INVX2 U7007 ( .A(DIN[8]), .Y(n6973) );
  INVX2 U7008 ( .A(DIN[7]), .Y(n6974) );
  INVX2 U7009 ( .A(DIN[6]), .Y(n6975) );
  INVX2 U7010 ( .A(DIN[5]), .Y(n6976) );
  INVX2 U7011 ( .A(DIN[4]), .Y(n6977) );
  INVX2 U7012 ( .A(DIN[3]), .Y(n6978) );
  INVX2 U7013 ( .A(DIN[31]), .Y(n6979) );
  INVX2 U7014 ( .A(DIN[30]), .Y(n6980) );
  INVX2 U7015 ( .A(DIN[2]), .Y(n6981) );
  INVX2 U7016 ( .A(DIN[29]), .Y(n6982) );
  INVX2 U7017 ( .A(DIN[28]), .Y(n6983) );
  INVX2 U7018 ( .A(DIN[27]), .Y(n6984) );
  INVX2 U7019 ( .A(DIN[26]), .Y(n6985) );
  INVX2 U7020 ( .A(DIN[25]), .Y(n6986) );
  INVX2 U7021 ( .A(DIN[24]), .Y(n6987) );
  INVX2 U7022 ( .A(DIN[23]), .Y(n6988) );
  INVX2 U7023 ( .A(DIN[22]), .Y(n6989) );
  INVX2 U7024 ( .A(DIN[21]), .Y(n6990) );
  INVX2 U7025 ( .A(DIN[20]), .Y(n6991) );
  INVX2 U7026 ( .A(DIN[1]), .Y(n6992) );
  INVX2 U7027 ( .A(DIN[19]), .Y(n6993) );
  INVX2 U7028 ( .A(DIN[18]), .Y(n6994) );
  INVX2 U7029 ( .A(DIN[17]), .Y(n6995) );
  INVX2 U7030 ( .A(DIN[16]), .Y(n6996) );
  INVX2 U7031 ( .A(DIN[15]), .Y(n6997) );
  INVX2 U7032 ( .A(DIN[14]), .Y(n6998) );
  INVX2 U7033 ( .A(DIN[13]), .Y(n6999) );
  INVX2 U7034 ( .A(DIN[12]), .Y(n7000) );
  INVX2 U7035 ( .A(DIN[11]), .Y(n7001) );
  INVX2 U7036 ( .A(DIN[10]), .Y(n7002) );
  INVX2 U7037 ( .A(DIN[0]), .Y(n7003) );
  INVX2 U7038 ( .A(n2217), .Y(n7004) );
  INVX2 U7039 ( .A(n889), .Y(n7005) );
  INVX2 U7040 ( .A(n622), .Y(n7006) );
  INVX2 U7041 ( .A(n354), .Y(n7007) );
  INVX2 U7042 ( .A(n1955), .Y(n7008) );
  INVX2 U7043 ( .A(n1688), .Y(n7009) );
  INVX2 U7044 ( .A(n1422), .Y(n7010) );
  INVX2 U7045 ( .A(n1155), .Y(n7011) );
  INVX2 U7046 ( .A(ADDR_WR[6]), .Y(n7012) );
  INVX2 U7047 ( .A(ADDR_WR[5]), .Y(n7013) );
  INVX2 U7048 ( .A(ADDR_WR[4]), .Y(n7014) );
  INVX2 U7049 ( .A(ADDR_WR[3]), .Y(n7015) );
  INVX2 U7050 ( .A(n2024), .Y(n7016) );
  INVX2 U7051 ( .A(n2061), .Y(n7017) );
  INVX2 U7052 ( .A(n2095), .Y(n7018) );
  INVX2 U7053 ( .A(n2129), .Y(n7019) );
  INVX2 U7054 ( .A(ADDR_WR[2]), .Y(n7020) );
  INVX2 U7055 ( .A(n1954), .Y(n7021) );
  INVX2 U7056 ( .A(n2163), .Y(n7022) );
  INVX2 U7057 ( .A(n2197), .Y(n7023) );
  INVX2 U7058 ( .A(n2220), .Y(n7024) );
  INVX2 U7059 ( .A(ADDR_WR[1]), .Y(n7025) );
  INVX2 U7060 ( .A(ADDR_WR[0]), .Y(n7026) );
endmodule


module ahb_slave ( clk, reset, HSEL, HADDR, HBURST, HSIZE, HTRANS, HWRITE, 
        HWDATA, RANDSPLIT, HMASTER, HMASTLOCK, HRDATA, HREADY, HRESP, HSPLIT, 
        STALL_pre );
  input [23:0] HADDR;
  input [2:0] HBURST;
  input [1:0] HSIZE;
  input [1:0] HTRANS;
  input [31:0] HWDATA;
  input [2:0] RANDSPLIT;
  input [3:0] HMASTER;
  output [31:0] HRDATA;
  output [1:0] HRESP;
  output [15:0] HSPLIT;
  input clk, reset, HSEL, HWRITE, HMASTLOCK, STALL_pre;
  output HREADY;
  wire   WR, RD;
  wire   [8:0] ADDR_WR;
  wire   [8:0] ADDR_RD;
  wire   [31:0] DIN;
  wire   [31:0] DOUT;

  ahb_slave_ram ahb_slave_ram ( .clk(clk), .reset(reset), .HSEL(HSEL), .HADDR(
        HADDR), .HBURST(HBURST), .HSIZE(HSIZE), .HTRANS(HTRANS), .HWRITE(
        HWRITE), .HWDATA(HWDATA), .RANDSPLIT(RANDSPLIT), .HMASTER(HMASTER), 
        .HMASTLOCK(HMASTLOCK), .HRDATA(HRDATA), .HREADY(HREADY), .HRESP(HRESP), 
        .HSPLIT(HSPLIT), .WR(WR), .RD(RD), .ADDR_WR(ADDR_WR), .ADDR_RD(ADDR_RD), .DIN(DIN), .DOUT(DOUT), .STALL_pre(STALL_pre) );
  ahb_slave_mem ahb_slave_mem ( .clk(clk), .reset(reset), .WR(WR), .RD(RD), 
        .ADDR_WR(ADDR_WR), .ADDR_RD(ADDR_RD), .DIN(DIN), .DOUT(DOUT) );
endmodule

